///////////////////////////////////////////////////////////////////////////////
//$Date: 2008/07/23 00:15:51 $
//$RCSfile: example_mgt_top.ejava,v $
//$Revision: 1.1.2.6 $
////////////////////////////////////////////////////////////////////////////////
//   ____  ____ 
//  /   /\/   / 
// /___/  \  /    Vendor: Xilinx 
// \   \   \/     Version : 1.5
//  \   \         Application : GTX Wizard 
//  /   /         Filename : example_mgt_top.v
// /___/   /\     Timestamp : 
// \   \  /  \ 
//  \___\/\___\ 
//
//
// Module EXAMPLE_MGT_TOP
// Generated by Xilinx GTX Wizard




`timescale 1ns / 1ps
`define DLY #1


//***********************************Entity Declaration************************

module EXAMPLE_MGT_TOP #
(
    parameter EXAMPLE_CONFIG_INDEPENDENT_LANES          =   1,   //configuration for frame gen and check
    parameter EXAMPLE_LANE_WITH_START_CHAR              =   0,   // specifies lane with unique start frame char
    parameter EXAMPLE_WORDS_IN_BRAM                     =   512, // specifies amount of data in BRAM 
    parameter EXAMPLE_SIM_MODE                          =   "FAST",  // Set to Fast Functional Simulation Model
    parameter EXAMPLE_SIM_GTXRESET_SPEEDUP              =   1,   // simulation setting for MGT smartmodel
    parameter EXAMPLE_SIM_PLL_PERDIV2                   =   9'h140, // simulation setting for MGT smartmodel
    parameter EXAMPLE_USE_CHIPSCOPE                     =   1    // Set to 1 to use Chipscope to drive resets
)
(
    TILE0_REFCLK_PAD_N_IN,
    TILE0_REFCLK_PAD_P_IN,
    GTXRESET_IN,
    TILE0_PLLLKDET_OUT,
    RXN_IN,
    RXP_IN,
    TXN_OUT,
    TXP_OUT
);

// synthesis attribute X_CORE_INFO of EXAMPLE_MGT_TOP is "gtxwizard_v1_5, Coregen v10.1_ip3";

//***********************************Ports Declaration*******************************

    input           TILE0_REFCLK_PAD_N_IN;
    input           TILE0_REFCLK_PAD_P_IN;
    input           GTXRESET_IN;
    output          TILE0_PLLLKDET_OUT;
    input   [1:0]   RXN_IN;
    input   [1:0]   RXP_IN;
    output  [1:0]   TXN_OUT;
    output  [1:0]   TXP_OUT;

    
//************************** Register Declarations ****************************

    reg     [84:0]  ila_in0_r;
    reg     [84:0]  ila_in1_r;
    reg             tile0_tx_resetdone1_r;
    reg             tile0_tx_resetdone1_r2;
    reg             tile0_rx_resetdone1_r;
    reg             tile0_rx_resetdone1_r2;
    

//**************************** Wire Declarations ******************************

    //------------------------ MGT Wrapper Wires ------------------------------
    

    //________________________________________________________________________
    //________________________________________________________________________
    //TILE0   (X0Y5)

    //---------------------- Loopback and Powerdown Ports ----------------------
    wire    [2:0]   tile0_loopback0_i;
    wire    [2:0]   tile0_loopback1_i;
    //--------------------- Receive Ports - 8b10b Decoder ----------------------
    wire            tile0_rxcharisk1_i;
    wire            tile0_rxdisperr1_i;
    wire            tile0_rxnotintable1_i;
    //----------------- Receive Ports - Clock Correction Ports -----------------
    wire    [2:0]   tile0_rxclkcorcnt1_i;
    //------------- Receive Ports - Comma Detection and Alignment --------------
    wire            tile0_rxenmcommaalign0_i;
    wire            tile0_rxenmcommaalign1_i;
    wire            tile0_rxenpcommaalign0_i;
    wire            tile0_rxenpcommaalign1_i;
    //----------------- Receive Ports - RX Data Path interface -----------------
    wire    [7:0]   tile0_rxdata1_i;
    wire            tile0_rxreset0_i;
    //------------- Receive Ports - RX Loss-of-sync State Machine --------------
    wire    [1:0]   tile0_rxlossofsync1_i;
    //------------------- Shared Ports - Tile and PLL Ports --------------------
    wire            tile0_gtxreset_i;
    wire            tile0_plllkdet_i;
    wire            tile0_refclkout_i;
    wire            tile0_resetdone0_i;
    wire            tile0_resetdone1_i;
    //-------------- Transmit Ports - 8b10b Encoder Control Ports --------------
    wire            tile0_txcharisk1_i;
    //---------------- Transmit Ports - TX Data Path interface -----------------
    wire    [7:0]   tile0_txdata1_i;


    //----------------------------- Global Signals -----------------------------
    wire            tile0_tx_system_reset0_c;
    wire            tile0_rx_system_reset0_c;
    wire            tile0_tx_system_reset1_c;
    wire            tile0_rx_system_reset1_c;
    wire            tied_to_ground_i;
    wire    [63:0]  tied_to_ground_vec_i;
    wire            tied_to_vcc_i;
    wire    [7:0]   tied_to_vcc_vec_i;
    wire            drp_clk_in_i;
    
    wire            tile0_refclkout_bufg_i;
    
    
    //--------------------------- User Clocks ---------------------------------
    wire            tile0_txusrclk1_i;
    wire            tile0_txusrclk21_i;
    wire            refclkout_pll0_locked_i;
    wire            refclkout_pll0_reset_i;
    wire            tile0_refclkout_to_cmt_i;


    //--------------------- Frame check/gen Module Signals --------------------
    wire            tile0_refclk_i;
    wire            tile0_matchn0_i;
    
    wire    [2:0]   tile0_txcharisk0_float_i;
    
    wire    [29:0]  tile0_txdata0_float_i;
    
    
    wire            tile0_block_sync0_reset_i;
    wire    [7:0]   tile0_error_count0_i;
    wire            tile0_frame_check0_reset_i;
    wire            tile0_inc_in0_i;
    wire            tile0_inc_out0_i;
    wire    [9:0]   tile0_unscrambled_data0_i;
    wire            tile0_matchn1_i;
    
    wire    [2:0]   tile0_txcharisk1_float_i;
    
    wire    [31:0]  tile0_txdata1_float_i;
    
    
    wire            tile0_block_sync1_reset_i;
    wire    [7:0]   tile0_error_count1_i;
    wire            tile0_frame_check1_reset_i;
    wire            tile0_inc_in1_i;
    wire            tile0_inc_out1_i;
    wire    [7:0]   tile0_unscrambled_data1_i;

    wire            reset_on_data_error_i;


    //--------------------- Chipscope Signals ---------------------------------

    wire    [35:0]  shared_vio_control_i;
    wire    [35:0]  tx_data_vio_control0_i;
    wire    [35:0]  tx_data_vio_control1_i;
    wire    [35:0]  rx_data_vio_control0_i;
    wire    [35:0]  rx_data_vio_control1_i;
    wire    [35:0]  ila_control0_i;
    wire    [35:0]  ila_control1_i;
    wire    [31:0]  shared_vio_in_i;
    wire    [31:0]  shared_vio_out_i;
    wire    [31:0]  tx_data_vio_in0_i;
    wire    [31:0]  tx_data_vio_out0_i;
    wire    [31:0]  tx_data_vio_in1_i;
    wire    [31:0]  tx_data_vio_out1_i;
    wire    [31:0]  rx_data_vio_in0_i;
    wire    [31:0]  rx_data_vio_out0_i;
    wire    [31:0]  rx_data_vio_in1_i;
    wire    [31:0]  rx_data_vio_out1_i;
    wire    [84:0]  ila_in0_i;
    wire    [84:0]  ila_in1_i;

    wire    [31:0]  tile0_tx_data_vio_in0_i;
    wire    [31:0]  tile0_tx_data_vio_out0_i;
    wire    [31:0]  tile0_tx_data_vio_in1_i;
    wire    [31:0]  tile0_tx_data_vio_out1_i;
    wire    [31:0]  tile0_rx_data_vio_in0_i;
    wire    [31:0]  tile0_rx_data_vio_out0_i;
    wire    [31:0]  tile0_rx_data_vio_in1_i;
    wire    [31:0]  tile0_rx_data_vio_out1_i;
    wire    [84:0]  tile0_ila_in0_i;
    wire    [84:0]  tile0_ila_in1_i;


    wire            gtxreset_i;
    wire            user_tx_reset_i;
    wire            user_rx_reset_i;
    wire            ila_clk0_i;
    wire            ila_clk_mux_out0_i;
    wire            ila_clk1_i;
    wire            ila_clk_mux_out1_i;


//**************************** Main Body of Code *******************************

    //  Static signal Assigments    
    assign tied_to_ground_i             = 1'b0;
    assign tied_to_ground_vec_i         = 64'h0000000000000000;
    assign tied_to_vcc_i                = 1'b1;
    assign tied_to_vcc_vec_i            = 8'hff;


    


    //---------------------Dedicated GTX Reference Clock Inputs ---------------
    // The dedicated reference clock inputs you selected in the GUI are implemented using
    // IBUFDS instances.
    //
    // In the UCF file for this example design, you will see that each of
    // these IBUFDS instances has been LOCed to a particular set of pins. By LOCing to these
    // locations, we tell the tools to use the dedicated input buffers to the GTX reference
    // clock network, rather than general purpose IOs. To select other pins, consult the 
    // Implementation chapter of UG196, or rerun the wizard.
    //
    // This network is the highest performace (lowest jitter) option for providing clocks
    // to the GTX transceivers.
    
    IBUFDS tile0_refclk_ibufds_i
    (
        .O                              (tile0_refclk_i), 
        .I                              (TILE0_REFCLK_PAD_P_IN),
        .IB                             (TILE0_REFCLK_PAD_N_IN)
    );






    //--------------------------------- User Clocks ---------------------------
    
    // The clock resources in this section were added based on userclk source selections on
    // the Latency, Buffering, and Clocking page of the GUI. A few notes about user clocks:
    // * The userclk and userclk2 for each GTX datapath (TX and RX) must be phase aligned to 
    //   avoid data errors in the fabric interface whenever the datapath is wider than 10 bits
    // * To minimize clock resources, you can share clocks between GTXs. GTXs using the same frequency
    //   or multiples of the same frequency can be accomadated using DCMs and PLLs. Use caution when
    //   using RXRECCLK as a clock source, however - these clocks can typically only be shared if all
    //   the channels using the clock are receiving data from TX channels that share a reference clock 
    //   source with each other.

    BUFG refclkout_pll0_bufg_i
    (
        .I                              (tile0_refclkout_i),
        .O                              (tile0_refclkout_to_cmt_i)
    );

    assign  refclkout_pll0_reset_i          =  !tile0_plllkdet_i;
    MGT_USRCLK_SOURCE_PLL #
    (
        .MULT                           (45),
        .DIVIDE                         (4),
        .CLK_PERIOD                     (16.0),
        .OUT0_DIVIDE                    (18),
        .OUT1_DIVIDE                    (9),
        .OUT2_DIVIDE                    (1),
        .OUT3_DIVIDE                    (1),
        .SIMULATION_P                   (EXAMPLE_USE_CHIPSCOPE),
        .LOCK_WAIT_COUNT                (16'b0001100001101010)
    )
    refclkout_pll0_i
    (
        .CLK0_OUT                       (tile0_txusrclk1_i),
        .CLK1_OUT                       (tile0_txusrclk21_i),
        .CLK2_OUT                       (),
        .CLK3_OUT                       (),
        .CLK_IN                         (tile0_refclkout_to_cmt_i),
        .PLL_LOCKED_OUT                 (refclkout_pll0_locked_i),
        .PLL_RESET_IN                   (refclkout_pll0_reset_i)
    );






    //--------------------------- The GTX Wrapper -----------------------------
    
    // Use the instantiation template in the examples directory to add the GTX wrapper to your design.
    // In this example, the wrapper is wired up for basic operation with a frame generator and frame 
    // checker. The GTXs will reset, then attempt to align and transmit data. If channel bonding is 
    // enabled, bonding should occur after alignment.
 
    // All clock inputs on the individual GTX transceiver must be driven for RESETDONE to work. 
    // When TX line Rate is set to No Tx, the source of TXUSRCLK(2) is set to rxusrclk(2).
    // When RX Line Rate is set to No RX, the source of RXUSRCLK(2) is set to txusrclk(2). 
    
    // Wire all PLLLKDET signals to the top level as output ports
    assign TILE0_PLLLKDET_OUT = tile0_plllkdet_i;


    ROCKETIO_GTX #
    (
        .WRAPPER_SIM_MODE               (EXAMPLE_SIM_MODE),
        .WRAPPER_SIM_GTXRESET_SPEEDUP   (EXAMPLE_SIM_GTXRESET_SPEEDUP),
        .WRAPPER_SIM_PLL_PERDIV2        (EXAMPLE_SIM_PLL_PERDIV2)
    )
    rocketio_gtx_i
    (
    
 
 
 
 
        //_____________________________________________________________________
        //_____________________________________________________________________
        //TILE0  (X0Y5)

        //---------------------- Loopback and Powerdown Ports ----------------------
        .TILE0_LOOPBACK0_IN             (tile0_loopback0_i),
        .TILE0_LOOPBACK1_IN             (tile0_loopback1_i),
        //--------------------- Receive Ports - 8b10b Decoder ----------------------
        .TILE0_RXCHARISK1_OUT           (tile0_rxcharisk1_i),
        .TILE0_RXDISPERR1_OUT           (tile0_rxdisperr1_i),
        .TILE0_RXNOTINTABLE1_OUT        (tile0_rxnotintable1_i),
        //----------------- Receive Ports - Clock Correction Ports -----------------
        .TILE0_RXCLKCORCNT1_OUT         (tile0_rxclkcorcnt1_i),
        //------------- Receive Ports - Comma Detection and Alignment --------------
        .TILE0_RXENMCOMMAALIGN0_IN      (tile0_rxenmcommaalign0_i),
        .TILE0_RXENMCOMMAALIGN1_IN      (tile0_rxenmcommaalign1_i),
        .TILE0_RXENPCOMMAALIGN0_IN      (tile0_rxenpcommaalign0_i),
        .TILE0_RXENPCOMMAALIGN1_IN      (tile0_rxenpcommaalign1_i),
        //----------------- Receive Ports - RX Data Path interface -----------------
        .TILE0_RXDATA1_OUT              (tile0_rxdata1_i),
        .TILE0_RXRESET0_IN              (tile0_rxreset0_i),
        .TILE0_RXRESET1_IN              (!refclkout_pll0_locked_i),
        .TILE0_RXUSRCLK0_IN             (tied_to_ground_i),
        .TILE0_RXUSRCLK1_IN             (tile0_txusrclk1_i),
        .TILE0_RXUSRCLK20_IN            (tied_to_ground_i),
        .TILE0_RXUSRCLK21_IN            (tile0_txusrclk21_i),
        //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        .TILE0_RXN0_IN                  (RXN_IN[0]),
        .TILE0_RXN1_IN                  (RXN_IN[1]),
        .TILE0_RXP0_IN                  (RXP_IN[0]),
        .TILE0_RXP1_IN                  (RXP_IN[1]),
        //------------- Receive Ports - RX Loss-of-sync State Machine --------------
        .TILE0_RXLOSSOFSYNC1_OUT        (tile0_rxlossofsync1_i),
        //------------------- Shared Ports - Tile and PLL Ports --------------------
        .TILE0_CLKIN_IN                 (tile0_refclk_i),
        .TILE0_GTXRESET_IN              (tile0_gtxreset_i),
        .TILE0_PLLLKDET_OUT             (tile0_plllkdet_i),
        .TILE0_REFCLKOUT_OUT            (tile0_refclkout_i),
        .TILE0_RESETDONE0_OUT           (tile0_resetdone0_i),
        .TILE0_RESETDONE1_OUT           (tile0_resetdone1_i),
        //-------------- Transmit Ports - 8b10b Encoder Control Ports --------------
        .TILE0_TXCHARISK1_IN            (tile0_txcharisk1_i),
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .TILE0_TXDATA1_IN               (tile0_txdata1_i),
        .TILE0_TXUSRCLK0_IN             (tied_to_ground_i),
        .TILE0_TXUSRCLK1_IN             (tile0_txusrclk1_i),
        .TILE0_TXUSRCLK20_IN            (tied_to_ground_i),
        .TILE0_TXUSRCLK21_IN            (tile0_txusrclk21_i),
        //------------- Transmit Ports - TX Driver and OOB signalling --------------
        .TILE0_TXN0_OUT                 (TXN_OUT[0]),
        .TILE0_TXN1_OUT                 (TXN_OUT[1]),
        .TILE0_TXP0_OUT                 (TXP_OUT[0]),
        .TILE0_TXP1_OUT                 (TXP_OUT[1])


    );







    //------------------------ User Module Resets -----------------------------
    // All the User Modules i.e. FRAME_GEN, FRAME_CHECK and the sync modules
    // are held in reset till the RESETDONE goes high. 
    // The RESETDONE is registered a couple of times on *USRCLK2 and connected 
    // to the reset of the modules
    
    
    always @(posedge tile0_txusrclk21_i or negedge tile0_resetdone1_i)

    begin
        if (!tile0_resetdone1_i )
        begin
            tile0_rx_resetdone1_r    <=   `DLY 1'b0;
            tile0_rx_resetdone1_r2   <=   `DLY 1'b0;
        end
        else
        begin
            tile0_rx_resetdone1_r    <=   `DLY tile0_resetdone1_i;
            tile0_rx_resetdone1_r2   <=   `DLY tile0_rx_resetdone1_r;
        end
    end
    
    
    always @(posedge tile0_txusrclk21_i or negedge tile0_resetdone1_i)

    begin
        if (!tile0_resetdone1_i )
        begin
            tile0_tx_resetdone1_r    <=   `DLY 1'b0;
            tile0_tx_resetdone1_r2   <=   `DLY 1'b0;
        end
        else
        begin
            tile0_tx_resetdone1_r    <=   `DLY tile0_resetdone1_i;
            tile0_tx_resetdone1_r2   <=   `DLY tile0_tx_resetdone1_r;
        end
    end

    



    //---------------------------- Frame Generators ---------------------------
    // The example design uses Block RAM based frame generators to provide test
    // data to the GTXs for transmission. By default the frame generators are 
    // loaded with an incrementing data sequence that includes commas/alignment
    // characters for alignment. If your protocol uses channel bonding, the 
    // frame generator will also be preloaded with a channel bonding sequence.
    
    // You can modify the data transmitted by changing the INIT values of the frame
    // generator in this file. Pay careful attention to bit order and the spacing
    // of your control and alignment characters.

    FRAME_GEN #
    (
        .WORDS_IN_BRAM(EXAMPLE_WORDS_IN_BRAM),
        .MEM_00(256'h0000000600000005000000040000000300000002000000bc0000000100000000),
        .MEM_01(256'h0000000e0000000d0000000c0000000b0000000a000000090000000800000007),
        .MEM_02(256'h000000160000001500000014000000130000001200000011000000100000000f),
        .MEM_03(256'h0000001e0000001d0000001c0000001b0000001a000000190000001800000017),
        .MEM_04(256'h000000260000002500000024000000230000002200000021000000200000001f),
        .MEM_05(256'h0000002e0000002d0000002c0000002b0000002a000000290000002800000027),
        .MEM_06(256'h000000360000003500000034000000330000003200000031000000300000002f),
        .MEM_07(256'h0000003e0000003d0000003c0000003b0000003a000000390000003800000037),
        .MEM_08(256'h000000460000004500000044000000430000004200000041000000400000003f),
        .MEM_09(256'h0000004e0000004d0000004c0000004b0000004a000000490000004800000047),
        .MEM_0A(256'h000000560000005500000054000000530000005200000051000000500000004f),
        .MEM_0B(256'h0000005e0000005d0000005c0000005b0000005a000000590000005800000057),
        .MEM_0C(256'h000000660000006500000064000000630000006200000061000000600000005f),
        .MEM_0D(256'h0000006e0000006d0000006c0000006b0000006a000000690000006800000067),
        .MEM_0E(256'h000000760000007500000074000000730000007200000071000000700000006f),
        .MEM_0F(256'h0000007e0000007d0000007c0000007b0000007a000000790000007800000077),
        .MEM_10(256'h0000000600000005000000040000000300000002000000bc0000000100000000),
        .MEM_11(256'h0000000e0000000d0000000c0000000b0000000a000000090000000800000007),
        .MEM_12(256'h000000160000001500000014000000130000001200000011000000100000000f),
        .MEM_13(256'h0000001e0000001d0000001c0000001b0000001a000000190000001800000017),
        .MEM_14(256'h000000260000002500000024000000230000002200000021000000200000001f),
        .MEM_15(256'h0000002e0000002d0000002c0000002b0000002a000000290000002800000027),
        .MEM_16(256'h000000360000003500000034000000330000003200000031000000300000002f),
        .MEM_17(256'h0000003e0000003d0000003c0000003b0000003a000000390000003800000037),
        .MEM_18(256'h000000460000004500000044000000430000004200000041000000400000003f),
        .MEM_19(256'h0000004e0000004d0000004c0000004b0000004a000000490000004800000047),
        .MEM_1A(256'h000000560000005500000054000000530000005200000051000000500000004f),
        .MEM_1B(256'h0000005e0000005d0000005c0000005b0000005a000000590000005800000057),
        .MEM_1C(256'h000000660000006500000064000000630000006200000061000000600000005f),
        .MEM_1D(256'h0000006e0000006d0000006c0000006b0000006a000000690000006800000067),
        .MEM_1E(256'h000000760000007500000074000000730000007200000071000000700000006f),
        .MEM_1F(256'h0000007e0000007d0000007c0000007b0000007a000000790000007800000077),
        .MEM_20(256'h0000000600000005000000040000000300000002000000bc0000000100000000),
        .MEM_21(256'h0000000e0000000d0000000c0000000b0000000a000000090000000800000007),
        .MEM_22(256'h000000160000001500000014000000130000001200000011000000100000000f),
        .MEM_23(256'h0000001e0000001d0000001c0000001b0000001a000000190000001800000017),
        .MEM_24(256'h000000260000002500000024000000230000002200000021000000200000001f),
        .MEM_25(256'h0000002e0000002d0000002c0000002b0000002a000000290000002800000027),
        .MEM_26(256'h000000360000003500000034000000330000003200000031000000300000002f),
        .MEM_27(256'h0000003e0000003d0000003c0000003b0000003a000000390000003800000037),
        .MEM_28(256'h000000460000004500000044000000430000004200000041000000400000003f),
        .MEM_29(256'h0000004e0000004d0000004c0000004b0000004a000000490000004800000047),
        .MEM_2A(256'h000000560000005500000054000000530000005200000051000000500000004f),
        .MEM_2B(256'h0000005e0000005d0000005c0000005b0000005a000000590000005800000057),
        .MEM_2C(256'h000000660000006500000064000000630000006200000061000000600000005f),
        .MEM_2D(256'h0000006e0000006d0000006c0000006b0000006a000000690000006800000067),
        .MEM_2E(256'h000000760000007500000074000000730000007200000071000000700000006f),
        .MEM_2F(256'h0000007e0000007d0000007c0000007b0000007a000000790000007800000077),
        .MEM_30(256'h0000000600000005000000040000000300000002000000bc0000000100000000),
        .MEM_31(256'h0000000e0000000d0000000c0000000b0000000a000000090000000800000007),
        .MEM_32(256'h000000160000001500000014000000130000001200000011000000100000000f),
        .MEM_33(256'h0000001e0000001d0000001c0000001b0000001a000000190000001800000017),
        .MEM_34(256'h000000260000002500000024000000230000002200000021000000200000001f),
        .MEM_35(256'h0000002e0000002d0000002c0000002b0000002a000000290000002800000027),
        .MEM_36(256'h000000360000003500000034000000330000003200000031000000300000002f),
        .MEM_37(256'h0000003e0000003d0000003c0000003b0000003a000000390000003800000037),
        .MEM_38(256'h000000460000004500000044000000430000004200000041000000400000003f),
        .MEM_39(256'h0000004e0000004d0000004c0000004b0000004a000000490000004800000047),
        .MEM_3A(256'h000000560000005500000054000000530000005200000051000000500000004f),
        .MEM_3B(256'h0000005e0000005d0000005c0000005b0000005a000000590000005800000057),
        .MEM_3C(256'h000000660000006500000064000000630000006200000061000000600000005f),
        .MEM_3D(256'h0000006e0000006d0000006c0000006b0000006a000000690000006800000067),
        .MEM_3E(256'h000000760000007500000074000000730000007200000071000000700000006f),
        .MEM_3F(256'h0000007e0000007d0000007c0000007b0000007a000000790000007800000077),
        .MEMP_00(256'h0000000000000000000000000000000000000000000000000000000000000100),
        .MEMP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .MEMP_02(256'h0000000000000000000000000000000000000000000000000000000000000100),
        .MEMP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .MEMP_04(256'h0000000000000000000000000000000000000000000000000000000000000100),
        .MEMP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .MEMP_06(256'h0000000000000000000000000000000000000000000000000000000000000100),
        .MEMP_07(256'h0000000000000000000000000000000000000000000000000000000000000000)
    )
    tile0_frame_gen1
    (
        // User Interface
        .TX_DATA                        ({tile0_txdata1_float_i,tile0_txdata1_i}),
    
    
        .TX_CHARISK                     ({tile0_txcharisk1_float_i,tile0_txcharisk1_i}),
    
        // System Interface
        .USER_CLK                       (tile0_txusrclk21_i),
        .SYSTEM_RESET                   (tile0_tx_system_reset1_c)
    );



    //-------------------------------- Frame Checkers -------------------------
    // The example design uses Block RAM based frame checkers to verify incoming  
    // data. By default the frame generators are loaded with a data sequence that 
    // matches the outgoing sequence of the frame generators for the TX ports.
    
    // You can modify the expected data sequence by changing the INIT values of the frame
    // checkers in this file. Pay careful attention to bit order and the spacing
    // of your control and alignment characters.
    
    // When the frame checker receives data, it attempts to synchronise to the 
    // incoming pattern by looking for the first sequence in the pattern. Once it 
    // finds the first sequence, it increments through the sequence, and indicates an 
    // error whenever the next value received does not match the expected value.

    
     // This GTX is not active.The match port for pattern checker of this GTX is tied off
     assign tile0_matchn0_i = 1'b0;


    assign tile0_frame_check1_reset_i = (EXAMPLE_CONFIG_INDEPENDENT_LANES==0)?reset_on_data_error_i:tile0_matchn1_i;

    // tile0_frame_check0 is always connected to the lane with the start of char
    // and this lane starts off the data checking on all the other lanes. The INC_IN port is tied off
    assign tile0_inc_in1_i = 1'b0;

    FRAME_CHECK #
    (
        .RX_DATA_WIDTH(8),
        .USE_COMMA(1),
        .WORDS_IN_BRAM(EXAMPLE_WORDS_IN_BRAM),
        .CONFIG_INDEPENDENT_LANES(1),
        .START_OF_PACKET_CHAR(8'hbc),
        .MEM_00(256'h0000000600000005000000040000000300000002000000bc0000000100000000),
        .MEM_01(256'h0000000e0000000d0000000c0000000b0000000a000000090000000800000007),
        .MEM_02(256'h000000160000001500000014000000130000001200000011000000100000000f),
        .MEM_03(256'h0000001e0000001d0000001c0000001b0000001a000000190000001800000017),
        .MEM_04(256'h000000260000002500000024000000230000002200000021000000200000001f),
        .MEM_05(256'h0000002e0000002d0000002c0000002b0000002a000000290000002800000027),
        .MEM_06(256'h000000360000003500000034000000330000003200000031000000300000002f),
        .MEM_07(256'h0000003e0000003d0000003c0000003b0000003a000000390000003800000037),
        .MEM_08(256'h000000460000004500000044000000430000004200000041000000400000003f),
        .MEM_09(256'h0000004e0000004d0000004c0000004b0000004a000000490000004800000047),
        .MEM_0A(256'h000000560000005500000054000000530000005200000051000000500000004f),
        .MEM_0B(256'h0000005e0000005d0000005c0000005b0000005a000000590000005800000057),
        .MEM_0C(256'h000000660000006500000064000000630000006200000061000000600000005f),
        .MEM_0D(256'h0000006e0000006d0000006c0000006b0000006a000000690000006800000067),
        .MEM_0E(256'h000000760000007500000074000000730000007200000071000000700000006f),
        .MEM_0F(256'h0000007e0000007d0000007c0000007b0000007a000000790000007800000077),
        .MEM_10(256'h0000000600000005000000040000000300000002000000bc0000000100000000),
        .MEM_11(256'h0000000e0000000d0000000c0000000b0000000a000000090000000800000007),
        .MEM_12(256'h000000160000001500000014000000130000001200000011000000100000000f),
        .MEM_13(256'h0000001e0000001d0000001c0000001b0000001a000000190000001800000017),
        .MEM_14(256'h000000260000002500000024000000230000002200000021000000200000001f),
        .MEM_15(256'h0000002e0000002d0000002c0000002b0000002a000000290000002800000027),
        .MEM_16(256'h000000360000003500000034000000330000003200000031000000300000002f),
        .MEM_17(256'h0000003e0000003d0000003c0000003b0000003a000000390000003800000037),
        .MEM_18(256'h000000460000004500000044000000430000004200000041000000400000003f),
        .MEM_19(256'h0000004e0000004d0000004c0000004b0000004a000000490000004800000047),
        .MEM_1A(256'h000000560000005500000054000000530000005200000051000000500000004f),
        .MEM_1B(256'h0000005e0000005d0000005c0000005b0000005a000000590000005800000057),
        .MEM_1C(256'h000000660000006500000064000000630000006200000061000000600000005f),
        .MEM_1D(256'h0000006e0000006d0000006c0000006b0000006a000000690000006800000067),
        .MEM_1E(256'h000000760000007500000074000000730000007200000071000000700000006f),
        .MEM_1F(256'h0000007e0000007d0000007c0000007b0000007a000000790000007800000077),
        .MEM_20(256'h0000000600000005000000040000000300000002000000bc0000000100000000),
        .MEM_21(256'h0000000e0000000d0000000c0000000b0000000a000000090000000800000007),
        .MEM_22(256'h000000160000001500000014000000130000001200000011000000100000000f),
        .MEM_23(256'h0000001e0000001d0000001c0000001b0000001a000000190000001800000017),
        .MEM_24(256'h000000260000002500000024000000230000002200000021000000200000001f),
        .MEM_25(256'h0000002e0000002d0000002c0000002b0000002a000000290000002800000027),
        .MEM_26(256'h000000360000003500000034000000330000003200000031000000300000002f),
        .MEM_27(256'h0000003e0000003d0000003c0000003b0000003a000000390000003800000037),
        .MEM_28(256'h000000460000004500000044000000430000004200000041000000400000003f),
        .MEM_29(256'h0000004e0000004d0000004c0000004b0000004a000000490000004800000047),
        .MEM_2A(256'h000000560000005500000054000000530000005200000051000000500000004f),
        .MEM_2B(256'h0000005e0000005d0000005c0000005b0000005a000000590000005800000057),
        .MEM_2C(256'h000000660000006500000064000000630000006200000061000000600000005f),
        .MEM_2D(256'h0000006e0000006d0000006c0000006b0000006a000000690000006800000067),
        .MEM_2E(256'h000000760000007500000074000000730000007200000071000000700000006f),
        .MEM_2F(256'h0000007e0000007d0000007c0000007b0000007a000000790000007800000077),
        .MEM_30(256'h0000000600000005000000040000000300000002000000bc0000000100000000),
        .MEM_31(256'h0000000e0000000d0000000c0000000b0000000a000000090000000800000007),
        .MEM_32(256'h000000160000001500000014000000130000001200000011000000100000000f),
        .MEM_33(256'h0000001e0000001d0000001c0000001b0000001a000000190000001800000017),
        .MEM_34(256'h000000260000002500000024000000230000002200000021000000200000001f),
        .MEM_35(256'h0000002e0000002d0000002c0000002b0000002a000000290000002800000027),
        .MEM_36(256'h000000360000003500000034000000330000003200000031000000300000002f),
        .MEM_37(256'h0000003e0000003d0000003c0000003b0000003a000000390000003800000037),
        .MEM_38(256'h000000460000004500000044000000430000004200000041000000400000003f),
        .MEM_39(256'h0000004e0000004d0000004c0000004b0000004a000000490000004800000047),
        .MEM_3A(256'h000000560000005500000054000000530000005200000051000000500000004f),
        .MEM_3B(256'h0000005e0000005d0000005c0000005b0000005a000000590000005800000057),
        .MEM_3C(256'h000000660000006500000064000000630000006200000061000000600000005f),
        .MEM_3D(256'h0000006e0000006d0000006c0000006b0000006a000000690000006800000067),
        .MEM_3E(256'h000000760000007500000074000000730000007200000071000000700000006f),
        .MEM_3F(256'h0000007e0000007d0000007c0000007b0000007a000000790000007800000077),
        .MEMP_00(256'h0000000000000000000000000000000000000000000000000000000000000100),
        .MEMP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .MEMP_02(256'h0000000000000000000000000000000000000000000000000000000000000100),
        .MEMP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .MEMP_04(256'h0000000000000000000000000000000000000000000000000000000000000100),
        .MEMP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .MEMP_06(256'h0000000000000000000000000000000000000000000000000000000000000100),
        .MEMP_07(256'h0000000000000000000000000000000000000000000000000000000000000000)
    )
    tile0_frame_check1
    (
        // MGT Interface
        .RX_DATA                        (tile0_rxdata1_i),  
        .RX_ENMCOMMA_ALIGN              (tile0_rxenmcommaalign1_i),
        .RX_ENPCOMMA_ALIGN              (tile0_rxenpcommaalign1_i),
        .RX_ENCHAN_SYNC                 ( ),
        .RX_CHANBOND_SEQ                (tied_to_ground_i),
        // Control Interface
        .INC_IN                         (tile0_inc_in1_i),
        .INC_OUT                        (tile0_inc_out1_i),
        .PATTERN_MATCH_N                (tile0_matchn1_i),
        .RESET_ON_ERROR                 (tile0_frame_check1_reset_i),
        // System Interface
        .USER_CLK                       (tile0_txusrclk21_i),
        .SYSTEM_RESET                   (tile0_rx_system_reset1_c),
        .ERROR_COUNT                    (tile0_error_count1_i)
  
    );

    





    //--------------------------- Chipscope Connections -----------------------
    // When the example design is run in hardware, it uses chipscope to allow the
    // example design and GTX wrapper to be controlled and monitored. The 
    // EXAMPLE_USE_CHIPSCOPE parameter allows chipscope to be removed for simulation.
    
generate
if (EXAMPLE_USE_CHIPSCOPE==1) 
begin : chipscope


    // Shared VIO for all tiles
    shared_vio shared_vio_i
    (
      .control                          (shared_vio_control_i),
      .async_in                         (shared_vio_in_i),
      .async_out                        (shared_vio_out_i)
    );

    // ICON for all VIOs 
    icon i_icon
    (
      .control0                         (shared_vio_control_i),
      .control1                         (tx_data_vio_control0_i),
      .control2                         (rx_data_vio_control0_i),
      .control3                         (ila_control0_i),
      .control4                         (tx_data_vio_control1_i),
      .control5                         (rx_data_vio_control1_i),
      .control6                         (ila_control1_i)
    );

    // TX VIO 
    shared_vio tx_data_vio0_i
    (
      .control                          (tx_data_vio_control0_i),
      .async_in                         (tx_data_vio_in0_i),
      .async_out                        (tx_data_vio_out0_i)  
    );
    
    // RX VIO 
    shared_vio rx_data_vio0_i
    (
      .control                          (rx_data_vio_control0_i),
      .async_in                         (rx_data_vio_in0_i),
      .async_out                        (rx_data_vio_out0_i)  
    );
    
    // RX ILA
    ila ila0_i
    (
      .control                          (ila_control0_i),
      .clk                              (ila_clk0_i),
      .trig0                            (ila_in0_i)
    );


    
    // The RX ILA must use the same clock as the selected transceiver
    BUFG ila_clk0_bufg_i
    (
        .I      (ila_clk_mux_out0_i),
        .O      (ila_clk0_i)
    );

    assign  ila_clk_mux_out0_i = 1'b0;


    // TX VIO 
    shared_vio tx_data_vio1_i
    (
      .control                          (tx_data_vio_control1_i),
      .async_in                         (tx_data_vio_in1_i),
      .async_out                        (tx_data_vio_out1_i)  
    );
    
    // RX VIO 
    shared_vio rx_data_vio1_i
    (
      .control                          (rx_data_vio_control1_i),
      .async_in                         (rx_data_vio_in1_i),
      .async_out                        (rx_data_vio_out1_i)  
    );
    
    // RX ILA
    ila ila1_i
    (
      .control                          (ila_control1_i),
      .clk                              (ila_clk1_i),
      .trig0                            (ila_in1_i)
    );


    
    // The RX ILA must use the same clock as the selected transceiver
    BUFG ila_clk1_bufg_i
    (
        .I      (ila_clk_mux_out1_i),
        .O      (ila_clk1_i)
    );

    assign  ila_clk_mux_out1_i = tile0_txusrclk21_i;



    // assign resets for frame_gen modules
    assign  tile0_tx_system_reset1_c = !tile0_tx_resetdone1_r2 || user_tx_reset_i;

    // assign resets for frame_check modules
    assign  tile0_rx_system_reset1_c = !tile0_rx_resetdone1_r2 || user_rx_reset_i;


    assign  tile0_gtxreset_i = gtxreset_i;

    // Shared VIO Outputs
    assign  gtxreset_i                      =  shared_vio_out_i[31];
    assign  user_tx_reset_i                 =  shared_vio_out_i[30];
    assign  user_rx_reset_i                 =  shared_vio_out_i[29];

    // Shared VIO Inputs
    assign  shared_vio_in_i[31]             =  tile0_plllkdet_i;
    assign  shared_vio_in_i[30:0]           =  31'b0000000000000000000000000000000;

    // Chipscope connections for GTP0 on Tile 0
    assign  tile0_tx_data_vio_in0_i[31:0]   =  32'b00000000000000000000000000000000;
    assign  tile0_loopback0_i               =  tx_data_vio_out0_i[31:29];
    assign  tile0_rx_data_vio_in0_i[31]     =  tile0_resetdone0_i;
    assign  tile0_rx_data_vio_in0_i[30:0]   =  31'b0000000000000000000000000000000;
    assign  tile0_ila_in0_i[84:77]          =  tile0_error_count0_i;
    assign  tile0_ila_in0_i[76:0]           =  77'b00000000000000000000000000000000000000000000000000000000000000000000000000000;

    // Chipscope connections for GTP1 on Tile 0
    assign  tile0_tx_data_vio_in1_i[31:0]   =  32'b00000000000000000000000000000000;
    assign  tile0_loopback1_i               =  tx_data_vio_out1_i[31:29];
    assign  tile0_rx_data_vio_in1_i[31]     =  tile0_resetdone1_i;
    assign  tile0_rx_data_vio_in1_i[30:0]   =  31'b0000000000000000000000000000000;
    assign  tile0_ila_in1_i[84]             =  tile0_rxcharisk1_i;
    assign  tile0_ila_in1_i[83]             =  tile0_rxdisperr1_i;
    assign  tile0_ila_in1_i[82]             =  tile0_rxnotintable1_i;
    assign  tile0_ila_in1_i[81:79]          =  tile0_rxclkcorcnt1_i;
    assign  tile0_ila_in1_i[78:71]          =  tile0_rxdata1_i;
    assign  tile0_ila_in1_i[70:69]          =  tile0_rxlossofsync1_i;
    assign  tile0_ila_in1_i[68:61]          =  tile0_error_count1_i;
    assign  tile0_ila_in1_i[60:0]           =  61'b0000000000000000000000000000000000000000000000000000000000000;



    assign  tx_data_vio_in0_i =                            tile0_tx_data_vio_in0_i;


    assign  rx_data_vio_in0_i =                            tile0_rx_data_vio_in0_i;


    assign  ila_in0_i =                                    tile0_ila_in0_i;


    assign  tx_data_vio_in1_i =                            tile0_tx_data_vio_in1_i;


    assign  rx_data_vio_in1_i =                            tile0_rx_data_vio_in1_i;


    assign  ila_in1_i =                                    tile0_ila_in1_i;




end //end EXAMPLE_USE_CHIPSCOPE=1 generate section
else 
begin: no_chipscope

    // If Chipscope is not being used, drive GTX reset signal
    // from the top level ports
    assign  tile0_gtxreset_i = GTXRESET_IN;

    // assign resets for frame_gen modules
    assign  tile0_tx_system_reset1_c = !tile0_tx_resetdone1_r2;

    // assign resets for frame_check modules
    assign  tile0_rx_system_reset1_c = !tile0_rx_resetdone1_r2;

    assign  gtxreset_i                      =  tied_to_ground_i;
    assign  user_tx_reset_i                 =  tied_to_ground_i;
    assign  user_rx_reset_i                 =  tied_to_ground_i;
    assign  tile0_loopback0_i               =  tied_to_ground_vec_i[2:0];
    assign  tile0_loopback1_i               =  tied_to_ground_vec_i[2:0];



end
endgenerate //End generate for EXAMPLE_USE_CHIPSCOPE


endmodule

//-------------------------------------------------------------------
//
//  VIO core module declaration 
//  This one is for driving shared ports and is asynchronous
//
//-------------------------------------------------------------------
module shared_vio
  (
    control,
    async_in,
    async_out
  );
  input  [35:0] control;
  input  [31:0] async_in;
  output [31:0] async_out;
endmodule

//-------------------------------------------------------------------
//
//  ICON core module declaration
//
//-------------------------------------------------------------------
module icon
  (
      control0,
      control1,
      control2,
      control3,
      control4,
      control5,
      control6  );
  output [35:0] control0;
  output [35:0] control1;
  output [35:0] control2;
  output [35:0] control3;
  output [35:0] control4;
  output [35:0] control5;
  output [35:0] control6;
endmodule


//-------------------------------------------------------------------
//
//  ILA core module declaration
//  This is used to allow RX signals to be monitored
//
//-------------------------------------------------------------------
module ila
  (
    control,
    clk,
    trig0
  );
  input [35:0] control;
  input clk;
  input [84:0] trig0;
endmodule


