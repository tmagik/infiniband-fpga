package ip_compatibility is
	type ip_provider_t is ( xilinx, altera );
end ip_compatibility;
