///////////////////////////////////////////////////////////////////////////////
//$Date: 2008/05/30 00:57:53 $
//$RCSfile: mgt_usrclk_source_dcm.ejava,v $
//$Revision: 1.1.2.1 $
///////////////////////////////////////////////////////////////////////////////
//   __  __ 
//  /   /\/   / 
// /__/  \   /    Vendor: Xilinx 
// \   \   \/     Version : 1.5
//  \   \         Application : RocketIO GTX Wizard 
//  /   /         Filename : mgt_usrclk_source.v
// /__/   /\      Timestamp : 02/08/2005 09:12:43
// \   \  /  \ 
//  \__\/\__\ 
//
//
// Module MGT_USRCLK_SOURCE (for use with GTX Transceivers)
// Generated by Xilinx RocketIO GTX Wizard

`timescale 1ns / 1ps

//***********************************Entity Declaration*******************************
module MGT_USRCLK_SOURCE #
(
    parameter FREQUENCY_MODE   = "LOW",
    parameter PERFORMANCE_MODE = "MAX_SPEED"
)
(
    DIV1_OUT,  
    DIV2_OUT,
    DCM_LOCKED_OUT,
    CLK_IN,  
    DCM_RESET_IN

);

// synthesis attribute X_CORE_INFO of MGT_USRCLK_SOURCE is "gtxwizard_v1_5, Coregen v10.1_ip3";

`define DLY #1


//*********************************** Port Declaration *******************************

    output          DIV1_OUT;
    output          DIV2_OUT;
    output          DCM_LOCKED_OUT;
    input           CLK_IN;
    input           DCM_RESET_IN;

//*********************************Wire Declarations**********************************

    wire    [15:0]  not_connected_i;
    wire            clkfb_i;
    wire            clkdv_i;
    wire            clk0_i;

//*********************************** Beginning of Code *******************************


    // Instantiate a DCM module to divide the reference clock.
    DCM_BASE #
    (
        .CLKDV_DIVIDE               (2.0),
        .DFS_FREQUENCY_MODE         ("LOW"), 
        .DLL_FREQUENCY_MODE         (FREQUENCY_MODE),    
        .DCM_PERFORMANCE_MODE       (PERFORMANCE_MODE)    
    )
    clock_divider_i
    (
        .CLK0                       (clk0_i),
        .CLK180                     (not_connected_i[0]),
        .CLK270                     (not_connected_i[1]),
        .CLK2X                      (not_connected_i[2]),
        .CLK2X180                   (not_connected_i[3]),
        .CLK90                      (not_connected_i[4]),
        .CLKDV                      (clkdv_i),
        .CLKFX                      (not_connected_i[5]),
        .CLKFX180                   (not_connected_i[6]),
        .LOCKED                     (DCM_LOCKED_OUT),
        .CLKFB                      (clkfb_i),
        .CLKIN                      (CLK_IN),
        .RST                        (DCM_RESET_IN)
    );

    
    BUFG dcm_1x_bufg_i
    (
        .I                          (clk0_i),
        .O                          (clkfb_i)
    );

    assign  DIV1_OUT  =   clkfb_i;


    BUFG dcm_div2_bufg_i
    (
        .I                          (clkdv_i),
        .O                          (DIV2_OUT)
    );


endmodule

