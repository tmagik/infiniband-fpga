------------------------------------------------------------------------------
--$Date: 2008/07/23 00:16:39 $
--$RCSfile: example_mgt_top_vhd.ejava,v $
--$Revision: 1.1.2.7 $
------------------------------------------------------------------------------
--   ____  ____ 
--  /   /\/   / 
-- /___/  \  /    Vendor: Xilinx 
-- \   \   \/     Version : 1.5
--  \   \         Application : RocketIO GTX Wizard 
--  /   /         Filename : example_mgt_top.vhd
-- /___/   /\     Timestamp : 
-- \   \  /  \ 
--  \___\/\___\ 
--
--
-- Module EXAMPLE_MGT_TOP
-- Generated by Xilinx RocketIO GTX Wizard

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;



--***********************************Entity Declaration************************

entity EXAMPLE_MGT_TOP is
generic
(
    EXAMPLE_CONFIG_INDEPENDENT_LANES        : integer   := 1;
    EXAMPLE_LANE_WITH_START_CHAR            : integer   := 0;
    EXAMPLE_WORDS_IN_BRAM                   : integer   := 512;
    EXAMPLE_SIM_MODE                        : string    := "FAST";
    EXAMPLE_SIM_GTXRESET_SPEEDUP            : integer   := 1;
    EXAMPLE_SIM_PLL_PERDIV2                 : bit_vector:= x"140";
    EXAMPLE_USE_CHIPSCOPE                   : integer   := 1     -- Set to 1 to use Chipscope to drive resets
);
port
(
    TILE0_REFCLK_PAD_N_IN                   : in   std_logic;
    TILE0_REFCLK_PAD_P_IN                   : in   std_logic;
    GTXRESET_IN                             : in   std_logic;
    TILE0_PLLLKDET_OUT                      : out  std_logic;
    RXN_IN                                  : in   std_logic_vector(1 downto 0);
    RXP_IN                                  : in   std_logic_vector(1 downto 0);
    TXN_OUT                                 : out  std_logic_vector(1 downto 0);
    TXP_OUT                                 : out  std_logic_vector(1 downto 0)
    
);

    attribute X_CORE_INFO : string;
    attribute X_CORE_INFO of EXAMPLE_MGT_TOP : entity is "gtxwizard_v1_5, Coregen v10.1_ip3";

end EXAMPLE_MGT_TOP;
    
architecture RTL of EXAMPLE_MGT_TOP is

--**************************Component Declarations*****************************


component ROCKETIO_GTX 
generic
(
    -- Simulation attributes
    WRAPPER_SIM_MODE                : string    := "FAST"; -- Set to Fast Functional Simulation Model
    WRAPPER_SIM_GTXRESET_SPEEDUP    : integer   := 0; -- Set to 1 to speed up sim reset
    WRAPPER_SIM_PLL_PERDIV2         : bit_vector:= x"140" -- Set to the VCO Unit Interval time
);
port
(
    
    --_________________________________________________________________________
    --_________________________________________________________________________
    --TILE0  (Location)

    ------------------------ Loopback and Powerdown Ports ----------------------
    TILE0_LOOPBACK0_IN                      : in   std_logic_vector(2 downto 0);
    TILE0_LOOPBACK1_IN                      : in   std_logic_vector(2 downto 0);
    ----------------------- Receive Ports - 8b10b Decoder ----------------------
    TILE0_RXCHARISK1_OUT                    : out  std_logic;
    TILE0_RXDISPERR1_OUT                    : out  std_logic;
    TILE0_RXNOTINTABLE1_OUT                 : out  std_logic;
    ------------------- Receive Ports - Clock Correction Ports -----------------
    TILE0_RXCLKCORCNT1_OUT                  : out  std_logic_vector(2 downto 0);
    --------------- Receive Ports - Comma Detection and Alignment --------------
    TILE0_RXENMCOMMAALIGN0_IN               : in   std_logic;
    TILE0_RXENMCOMMAALIGN1_IN               : in   std_logic;
    TILE0_RXENPCOMMAALIGN0_IN               : in   std_logic;
    TILE0_RXENPCOMMAALIGN1_IN               : in   std_logic;
    ------------------- Receive Ports - RX Data Path interface -----------------
    TILE0_RXDATA1_OUT                       : out  std_logic_vector(7 downto 0);
    TILE0_RXRESET0_IN                       : in   std_logic;
    TILE0_RXRESET1_IN                       : in   std_logic;
    TILE0_RXUSRCLK0_IN                      : in   std_logic;
    TILE0_RXUSRCLK1_IN                      : in   std_logic;
    TILE0_RXUSRCLK20_IN                     : in   std_logic;
    TILE0_RXUSRCLK21_IN                     : in   std_logic;
    ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    TILE0_RXN0_IN                           : in   std_logic;
    TILE0_RXN1_IN                           : in   std_logic;
    TILE0_RXP0_IN                           : in   std_logic;
    TILE0_RXP1_IN                           : in   std_logic;
    --------------- Receive Ports - RX Loss-of-sync State Machine --------------
    TILE0_RXLOSSOFSYNC1_OUT                 : out  std_logic_vector(1 downto 0);
    --------------------- Shared Ports - Tile and PLL Ports --------------------
    TILE0_CLKIN_IN                          : in   std_logic;
    TILE0_GTXRESET_IN                       : in   std_logic;
    TILE0_PLLLKDET_OUT                      : out  std_logic;
    TILE0_REFCLKOUT_OUT                     : out  std_logic;
    TILE0_RESETDONE0_OUT                    : out  std_logic;
    TILE0_RESETDONE1_OUT                    : out  std_logic;
    ---------------- Transmit Ports - 8b10b Encoder Control Ports --------------
    TILE0_TXCHARISK1_IN                     : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    TILE0_TXDATA1_IN                        : in   std_logic_vector(7 downto 0);
    TILE0_TXUSRCLK0_IN                      : in   std_logic;
    TILE0_TXUSRCLK1_IN                      : in   std_logic;
    TILE0_TXUSRCLK20_IN                     : in   std_logic;
    TILE0_TXUSRCLK21_IN                     : in   std_logic;
    --------------- Transmit Ports - TX Driver and OOB signalling --------------
    TILE0_TXN0_OUT                          : out  std_logic;
    TILE0_TXN1_OUT                          : out  std_logic;
    TILE0_TXP0_OUT                          : out  std_logic;
    TILE0_TXP1_OUT                          : out  std_logic


);
end component;


component MGT_USRCLK_SOURCE 
generic
(
    FREQUENCY_MODE   : string   := "LOW";    
    PERFORMANCE_MODE : string   := "MAX_SPEED"    
);
port
(
    DIV1_OUT                : out std_logic;
    DIV2_OUT                : out std_logic;
    DCM_LOCKED_OUT          : out std_logic;
    CLK_IN                  : in  std_logic;
    DCM_RESET_IN            : in  std_logic

);
end component;

component FRAME_GEN 
generic
(
    WORDS_IN_BRAM : integer    :=   256;
    MEM_00       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_01       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_02       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_03       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_04       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_05       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_06       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_07       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_08       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_09       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0A       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0B       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0C       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0D       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0E       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0F       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_10       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_11       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_12       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_13       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_14       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_15       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_16       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_17       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_18       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_19       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1A       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1B       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1C       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1D       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1E       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1F       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_20       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_21       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_22       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_23       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_24       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_25       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_26       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_27       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_28       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_29       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2A       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2B       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2C       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2D       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2E       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2F       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_30       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_31       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_32       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_33       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_34       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_35       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_36       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_37       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_38       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_39       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3A       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3B       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3C       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3D       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3E       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3F       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_00      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_01      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_02      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_03      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_04      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_05      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_06      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_07      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000"
);    
port
(
    -- User Interface
    TX_DATA             : out   std_logic_vector(39 downto 0);
    TX_CHARISK          : out   std_logic_vector(3 downto 0); 

    -- System Interface
    USER_CLK            : in    std_logic;
    SYSTEM_RESET        : in    std_logic
); 
end component;

component FRAME_CHECK 
generic
(
    RX_DATA_WIDTH            : integer := 16;
    USE_COMMA                : integer := 1;
    NONE_MSB_FIRST_DEC       : integer := 0;
    COMMA_DOUBLE_DEC         : integer := 0;
    CHANBOND_SEQ_LEN         : integer := 1;
    WORDS_IN_BRAM            : integer := 256;
    CONFIG_INDEPENDENT_LANES : integer := 0;
    START_OF_PACKET_CHAR     : std_logic_vector := x"55fb";
    COMMA_DOUBLE_CHAR        : std_logic_vector := x"f628";
    MEM_00       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_01       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_02       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_03       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_04       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_05       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_06       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_07       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_08       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_09       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0A       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0B       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0C       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0D       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0E       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0F       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_10       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_11       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_12       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_13       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_14       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_15       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_16       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_17       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_18       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_19       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1A       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1B       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1C       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1D       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1E       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1F       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_20       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_21       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_22       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_23       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_24       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_25       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_26       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_27       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_28       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_29       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2A       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2B       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2C       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2D       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2E       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2F       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_30       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_31       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_32       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_33       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_34       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_35       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_36       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_37       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_38       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_39       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3A       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3B       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3C       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3D       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3E       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3F       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_00      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_01      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_02      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_03      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_04      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_05      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_06      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_07      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000"
);
port
(
    -- User Interface
    RX_DATA                  : in  std_logic_vector((RX_DATA_WIDTH-1) downto 0); 
    RX_ENMCOMMA_ALIGN        : out std_logic;
    RX_ENPCOMMA_ALIGN        : out std_logic;
    RX_ENCHAN_SYNC           : out std_logic; 
    RX_CHANBOND_SEQ          : in  std_logic; 

    -- Control Interface
    INC_IN                   : in std_logic; 
    INC_OUT                  : out std_logic; 
    PATTERN_MATCH_N          : out std_logic;
    RESET_ON_ERROR           : in std_logic; 
    
    -- Error Monitoring
    ERROR_COUNT              : out std_logic_vector(7 downto 0);

    -- System Interface
    USER_CLK                 : in std_logic;
    SYSTEM_RESET             : in std_logic
  
);
end component;

component MGT_USRCLK_SOURCE_PLL 
generic
(
    MULT                 : integer          := 2;
    DIVIDE               : integer          := 2;    
    CLK_PERIOD           : real             := 16.0;    
    OUT0_DIVIDE          : integer          := 2;
    OUT1_DIVIDE          : integer          := 2;
    OUT2_DIVIDE          : integer          := 2;
    OUT3_DIVIDE          : integer          := 2;
    SIMULATION_P         : integer          := 1;
    LOCK_WAIT_COUNT      : std_logic_vector := "1000001000110101"  
);
port
( 
    CLK0_OUT                : out std_logic;
    CLK1_OUT                : out std_logic;
    CLK2_OUT                : out std_logic;
    CLK3_OUT                : out std_logic;
    CLK_IN                  : in  std_logic;
    PLL_LOCKED_OUT          : out std_logic;
    PLL_RESET_IN            : in  std_logic
);
end component;






-- Chipscope modules
attribute syn_black_box                : boolean;
attribute syn_noprune                  : boolean;


component shared_vio
port
(
    control                 : in  std_logic_vector(35 downto 0);
    async_in                : in  std_logic_vector(31 downto 0);
    async_out               : out std_logic_vector(31 downto 0)
);
end component;
attribute syn_black_box of shared_vio : component is TRUE;
attribute syn_noprune of shared_vio   : component is TRUE;

component icon
port
(
    control0                : out std_logic_vector(35 downto 0);
    control1                : out std_logic_vector(35 downto 0);
    control2                : out std_logic_vector(35 downto 0);
    control3                : out std_logic_vector(35 downto 0);
    control4                : out std_logic_vector(35 downto 0);
    control5                : out std_logic_vector(35 downto 0);
    control6                : out std_logic_vector(35 downto 0));
end component;


attribute syn_black_box of icon : component is TRUE;
attribute syn_noprune of icon   : component is TRUE;


component ila
port
(
    control                 : in  std_logic_vector(35 downto 0);
    clk                     : in  std_logic;
    trig0                   : in  std_logic_vector(84 downto 0)
);
end component;
attribute syn_black_box of ila : component is TRUE;
attribute syn_noprune of ila   : component is TRUE;


--***********************************Parameter Declarations********************

    constant DLY : time := 1 ns;

    
--************************** Register Declarations ****************************

    signal   tile0_tx_resetdone1_r           : std_logic;
    signal   tile0_tx_resetdone1_r2          : std_logic;
    signal   tile0_rx_resetdone1_r           : std_logic;
    signal   tile0_rx_resetdone1_r2          : std_logic;
  

--**************************** Wire Declarations ******************************

    -------------------------- MGT Wrapper Wires ------------------------------
    
    --________________________________________________________________________
    --________________________________________________________________________
    --TILE0   (X0Y5)

    ------------------------ Loopback and Powerdown Ports ----------------------
    signal  tile0_loopback0_i               : std_logic_vector(2 downto 0);
    signal  tile0_loopback1_i               : std_logic_vector(2 downto 0);
    ----------------------- Receive Ports - 8b10b Decoder ----------------------
    signal  tile0_rxcharisk1_i              : std_logic;
    signal  tile0_rxdisperr1_i              : std_logic;
    signal  tile0_rxnotintable1_i           : std_logic;
    ------------------- Receive Ports - Clock Correction Ports -----------------
    signal  tile0_rxclkcorcnt1_i            : std_logic_vector(2 downto 0);
    --------------- Receive Ports - Comma Detection and Alignment --------------
    signal  tile0_rxenmcommaalign0_i        : std_logic;
    signal  tile0_rxenmcommaalign1_i        : std_logic;
    signal  tile0_rxenpcommaalign0_i        : std_logic;
    signal  tile0_rxenpcommaalign1_i        : std_logic;
    ------------------- Receive Ports - RX Data Path interface -----------------
    signal  tile0_rxdata1_i                 : std_logic_vector(7 downto 0);
    signal  tile0_rxreset0_i                : std_logic;
    signal  tile0_rxreset1_i                : std_logic;
    --------------- Receive Ports - RX Loss-of-sync State Machine --------------
    signal  tile0_rxlossofsync1_i           : std_logic_vector(1 downto 0);
    --------------------- Shared Ports - Tile and PLL Ports --------------------
    signal  tile0_gtxreset_i                : std_logic;
    signal  tile0_plllkdet_i                : std_logic;
    signal  tile0_refclkout_i               : std_logic;
    signal  tile0_resetdone0_i              : std_logic;
    signal  tile0_resetdone1_i              : std_logic;
    ---------------- Transmit Ports - 8b10b Encoder Control Ports --------------
    signal  tile0_txcharisk1_i              : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  tile0_txdata1_i                 : std_logic_vector(7 downto 0);


    ------------------------------- Global Signals -----------------------------
    signal  tile0_tx_system_reset0_c        : std_logic;
    signal  tile0_rx_system_reset0_c        : std_logic;
    signal  tile0_tx_system_reset1_c        : std_logic;
    signal  tile0_rx_system_reset1_c        : std_logic;
    signal  tied_to_ground_i                : std_logic;
    signal  tied_to_ground_vec_i            : std_logic_vector(63 downto 0);
    signal  tied_to_vcc_i                   : std_logic;
    signal  tied_to_vcc_vec_i               : std_logic_vector(7 downto 0);
    signal  drp_clk_in_i                    : std_logic;
    
    signal  tile0_refclkout_bufg_i          : std_logic;
    
    
    ----------------------------- User Clocks ---------------------------------
    signal  tile0_txusrclk1_i               : std_logic;
    signal  tile0_txusrclk21_i              : std_logic;
    signal  refclkout_pll0_locked_i         : std_logic;
    signal  refclkout_pll0_reset_i          : std_logic;
    signal  tile0_refclkout_to_cmt_i        : std_logic;


    ----------------------- Frame check/gen Module Signals --------------------
    signal  tile0_refclk_i                  : std_logic;
    signal  tile0_matchn0_i                 : std_logic;
     
    signal  tile0_txcharisk0_float_i        : std_logic_vector(2 downto 0);
    signal  tile0_txdata0_float_i           : std_logic_vector(29 downto 0);
    
    
    signal  tile0_block_sync0_i             : std_logic;
    signal  tile0_error_count0_i            : std_logic_vector(7 downto 0);
    signal  tile0_frame_check0_reset_i      : std_logic;
    signal  tile0_inc_in0_i                 : std_logic;
    signal  tile0_inc_out0_i                : std_logic;
    signal  tile0_unscrambled_data0_i       : std_logic_vector(9 downto 0);
    signal  tile0_matchn1_i                 : std_logic;
     
    signal  tile0_txcharisk1_float_i        : std_logic_vector(2 downto 0);
    signal  tile0_txdata1_float_i           : std_logic_vector(31 downto 0);
    
    
    signal  tile0_block_sync1_i             : std_logic;
    signal  tile0_error_count1_i            : std_logic_vector(7 downto 0);
    signal  tile0_frame_check1_reset_i      : std_logic;
    signal  tile0_inc_in1_i                 : std_logic;
    signal  tile0_inc_out1_i                : std_logic;
    signal  tile0_unscrambled_data1_i       : std_logic_vector(7 downto 0);

    signal  reset_on_data_error_i           : std_logic;


    ----------------------- Chipscope Signals ---------------------------------

    signal  shared_vio_control_i            : std_logic_vector(35 downto 0);
    signal  tx_data_vio_control0_i          : std_logic_vector(35 downto 0);
    signal  tx_data_vio_control1_i          : std_logic_vector(35 downto 0);
    signal  rx_data_vio_control0_i          : std_logic_vector(35 downto 0);
    signal  rx_data_vio_control1_i          : std_logic_vector(35 downto 0);
    signal  ila_control0_i                  : std_logic_vector(35 downto 0);
    signal  ila_control1_i                  : std_logic_vector(35 downto 0);
    signal  shared_vio_in_i                 : std_logic_vector(31 downto 0);
    signal  shared_vio_out_i                : std_logic_vector(31 downto 0);
    signal  tx_data_vio_in0_i               : std_logic_vector(31 downto 0);
    signal  tx_data_vio_out0_i              : std_logic_vector(31 downto 0);
    signal  tx_data_vio_in1_i               : std_logic_vector(31 downto 0);
    signal  tx_data_vio_out1_i              : std_logic_vector(31 downto 0);
    signal  rx_data_vio_in0_i               : std_logic_vector(31 downto 0);
    signal  rx_data_vio_out0_i              : std_logic_vector(31 downto 0);
    signal  rx_data_vio_in1_i               : std_logic_vector(31 downto 0);
    signal  rx_data_vio_out1_i              : std_logic_vector(31 downto 0);
    signal  ila_in0_i                       : std_logic_vector(84 downto 0);
    signal  ila_in1_i                       : std_logic_vector(84 downto 0);

    signal  tile0_tx_data_vio_in0_i         : std_logic_vector(31 downto 0);
    signal  tile0_tx_data_vio_out0_i        : std_logic_vector(31 downto 0);
    signal  tile0_tx_data_vio_in1_i         : std_logic_vector(31 downto 0);
    signal  tile0_tx_data_vio_out1_i        : std_logic_vector(31 downto 0);
    signal  tile0_rx_data_vio_in0_i         : std_logic_vector(31 downto 0);
    signal  tile0_rx_data_vio_out0_i        : std_logic_vector(31 downto 0);
    signal  tile0_rx_data_vio_in1_i         : std_logic_vector(31 downto 0);
    signal  tile0_rx_data_vio_out1_i        : std_logic_vector(31 downto 0);
    signal  tile0_ila_in0_i                 : std_logic_vector(84 downto 0);
    signal  tile0_ila_in1_i                 : std_logic_vector(84 downto 0);


    signal  gtxreset_i                      : std_logic;
    signal  user_tx_reset_i                 : std_logic;
    signal  user_rx_reset_i                 : std_logic;
    signal  ila_clk0_i                      : std_logic;
    signal  ila_clk_mux_out0_i              : std_logic;
    signal  ila_clk1_i                      : std_logic;
    signal  ila_clk_mux_out1_i              : std_logic;


--**************************** Main Body of Code *******************************
begin

    --  Static signal Assigments
    tied_to_ground_i                        <= '0';
    tied_to_ground_vec_i                    <= x"0000000000000000";
    tied_to_vcc_i                           <= '1';
    tied_to_vcc_vec_i                       <= x"ff";


    


    -----------------------Dedicated GTX Reference Clock Inputs ---------------
    -- The dedicated reference clock inputs you selected in the GUI are implemented using
    -- IBUFDS instances.
    --
    -- In the UCF file for this example design, you will see that each of
    -- these IBUFDS instances has been LOCed to a particular set of pins. By LOCing to these
    -- locations, we tell the tools to use the dedicated input buffers to the GTX reference
    -- clock network, rather than general purpose IOs. To select other pins, consult the 
    -- Implementation chapter of UG196, or rerun the wizard.
    --
    -- This network is the highest performace (lowest jitter) option for providing clocks
    -- to the GTX transceivers.
    
    tile0_refclk_ibufds_i : IBUFDS
    port map
    (
        O                               =>      tile0_refclk_i,
        I                               =>      TILE0_REFCLK_PAD_P_IN,
        IB                              =>      TILE0_REFCLK_PAD_N_IN
    );






    ----------------------------------- User Clocks ---------------------------
    
    -- The clock resources in this section were added based on userclk source selections on
    -- the Latency, Buffering, and Clocking page of the GUI. A few notes about user clocks:
    -- * The userclk and userclk2 for each GTX datapath (TX and RX) must be phase aligned to 
    --   avoid data errors in the fabric interface whenever the datapath is wider than 10 bits
    -- * To minimize clock resources, you can share clocks between GTXs. GTXs using the same frequency
    --   or multiples of the same frequency can be accomadated using DCMs and PLLs. Use caution when
    --   using RXRECCLK as a clock source, however - these clocks can typically only be shared if all
    --   the channels using the clock are receiving data from TX channels that share a reference clock 
    --   source with each other.

    refclkout_pll0_bufg_i : BUFG
    port map
    (
        I                               =>      tile0_refclkout_i,
        O                               =>      tile0_refclkout_to_cmt_i
    );

    refclkout_pll0_reset_i                  <= not tile0_plllkdet_i;
    refclkout_pll0_i : MGT_USRCLK_SOURCE_PLL
    generic map
    (
        MULT                            =>      45,
        DIVIDE                          =>      4,
        CLK_PERIOD                      =>      16.0,
        OUT0_DIVIDE                     =>      18,
        OUT1_DIVIDE                     =>      9,
        OUT2_DIVIDE                     =>      1,
        OUT3_DIVIDE                     =>      1,
        SIMULATION_P                    =>      EXAMPLE_USE_CHIPSCOPE,
        LOCK_WAIT_COUNT                 =>      "0001100001101010"
    )
    port map
    (
        CLK0_OUT                        =>      tile0_txusrclk1_i,
        CLK1_OUT                        =>      tile0_txusrclk21_i,
        CLK2_OUT                        =>      open,
        CLK3_OUT                        =>      open,
        CLK_IN                          =>      tile0_refclkout_to_cmt_i,
        PLL_LOCKED_OUT                  =>      refclkout_pll0_locked_i,
        PLL_RESET_IN                    =>      refclkout_pll0_reset_i
    );






    ----------------------------- The GTX Wrapper -----------------------------
    
    -- Use the instantiation template in the examples directory to add the GTX wrapper to your design.
    -- In this example, the wrapper is wired up for basic operation with a frame generator and frame 
    -- checker. The GTXs will reset, then attempt to align and transmit data. If channel bonding is 
    -- enabled, bonding should occur after alignment.

    -- All clock inputs on the individual GTX transceiver must be driven for RESETDONE to work.
    -- When TX line Rate is set to No Tx, the source of TXUSRCLK(2) is set to rxusrclk(2).
    -- When RX Line Rate is set to No RX, the source of RXUSRCLK(2) is set to txusrclk(2). 

    -- Wire all PLLLKDET signals to the top level as output ports
    TILE0_PLLLKDET_OUT                      <= tile0_plllkdet_i;


    -- Hold the RX in reset till the RX user clocks are stable
  
    tile0_rxreset1_i                    <= not refclkout_pll0_locked_i;

    rocketio_gtx_i : ROCKETIO_GTX
    generic map
    (
        WRAPPER_SIM_MODE                =>      EXAMPLE_SIM_MODE,
        WRAPPER_SIM_GTXRESET_SPEEDUP    =>      EXAMPLE_SIM_GTXRESET_SPEEDUP,
        WRAPPER_SIM_PLL_PERDIV2         =>      EXAMPLE_SIM_PLL_PERDIV2
    )
    port map
    (
    
 
 
 
 
        --_____________________________________________________________________
        --_____________________________________________________________________
        --TILE0  (X0Y5)

        ------------------------ Loopback and Powerdown Ports ----------------------
        TILE0_LOOPBACK0_IN              =>      tile0_loopback0_i,
        TILE0_LOOPBACK1_IN              =>      tile0_loopback1_i,
        ----------------------- Receive Ports - 8b10b Decoder ----------------------
        TILE0_RXCHARISK1_OUT            =>      tile0_rxcharisk1_i,
        TILE0_RXDISPERR1_OUT            =>      tile0_rxdisperr1_i,
        TILE0_RXNOTINTABLE1_OUT         =>      tile0_rxnotintable1_i,
        ------------------- Receive Ports - Clock Correction Ports -----------------
        TILE0_RXCLKCORCNT1_OUT          =>      tile0_rxclkcorcnt1_i,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        TILE0_RXENMCOMMAALIGN0_IN       =>      tile0_rxenmcommaalign0_i,
        TILE0_RXENMCOMMAALIGN1_IN       =>      tile0_rxenmcommaalign1_i,
        TILE0_RXENPCOMMAALIGN0_IN       =>      tile0_rxenpcommaalign0_i,
        TILE0_RXENPCOMMAALIGN1_IN       =>      tile0_rxenpcommaalign1_i,
        ------------------- Receive Ports - RX Data Path interface -----------------
        TILE0_RXDATA1_OUT               =>      tile0_rxdata1_i,
        TILE0_RXRESET0_IN               =>      tile0_rxreset0_i,
        TILE0_RXRESET1_IN               =>      tile0_rxreset1_i,
        TILE0_RXUSRCLK0_IN              =>      tied_to_ground_i,
        TILE0_RXUSRCLK1_IN              =>      tile0_txusrclk1_i,
        TILE0_RXUSRCLK20_IN             =>      tied_to_ground_i,
        TILE0_RXUSRCLK21_IN             =>      tile0_txusrclk21_i,
        ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        TILE0_RXN0_IN                   =>      RXN_IN(0),
        TILE0_RXN1_IN                   =>      RXN_IN(1),
        TILE0_RXP0_IN                   =>      RXP_IN(0),
        TILE0_RXP1_IN                   =>      RXP_IN(1),
        --------------- Receive Ports - RX Loss-of-sync State Machine --------------
        TILE0_RXLOSSOFSYNC1_OUT         =>      tile0_rxlossofsync1_i,
        --------------------- Shared Ports - Tile and PLL Ports --------------------
        TILE0_CLKIN_IN                  =>      tile0_refclk_i,
        TILE0_GTXRESET_IN               =>      tile0_gtxreset_i,
        TILE0_PLLLKDET_OUT              =>      tile0_plllkdet_i,
        TILE0_REFCLKOUT_OUT             =>      tile0_refclkout_i,
        TILE0_RESETDONE0_OUT            =>      tile0_resetdone0_i,
        TILE0_RESETDONE1_OUT            =>      tile0_resetdone1_i,
        ---------------- Transmit Ports - 8b10b Encoder Control Ports --------------
        TILE0_TXCHARISK1_IN             =>      tile0_txcharisk1_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        TILE0_TXDATA1_IN                =>      tile0_txdata1_i,
        TILE0_TXUSRCLK0_IN              =>      tied_to_ground_i,
        TILE0_TXUSRCLK1_IN              =>      tile0_txusrclk1_i,
        TILE0_TXUSRCLK20_IN             =>      tied_to_ground_i,
        TILE0_TXUSRCLK21_IN             =>      tile0_txusrclk21_i,
        --------------- Transmit Ports - TX Driver and OOB signalling --------------
        TILE0_TXN0_OUT                  =>      TXN_OUT(0),
        TILE0_TXN1_OUT                  =>      TXN_OUT(1),
        TILE0_TXP0_OUT                  =>      TXP_OUT(0),
        TILE0_TXP1_OUT                  =>      TXP_OUT(1)


    );







    -------------------------- User Module Resets -----------------------------
    -- All the User Modules i.e. FRAME_GEN, FRAME_CHECK and the sync modules
    -- are held in reset till the RESETDONE goes high. 
    -- The RESETDONE is registered a couple of times on USRCLK2 and connected 
    -- to the reset of the modules
    
    process( tile0_txusrclk21_i,tile0_resetdone1_i)
    begin
        if(tile0_resetdone1_i = '0') then
            tile0_rx_resetdone1_r  <= '0'   after DLY;
            tile0_rx_resetdone1_r2 <= '0'   after DLY;
        elsif(tile0_txusrclk21_i'event and tile0_txusrclk21_i = '1') then
            tile0_rx_resetdone1_r  <= tile0_resetdone1_i   after DLY;
            tile0_rx_resetdone1_r2 <= tile0_rx_resetdone1_r   after DLY;
        end if;
    end process;
    process( tile0_txusrclk21_i,tile0_resetdone1_i)
    begin
        if(tile0_resetdone1_i = '0') then
            tile0_tx_resetdone1_r  <= '0'   after DLY;
            tile0_tx_resetdone1_r2 <= '0'   after DLY;
        elsif(tile0_txusrclk21_i'event and tile0_txusrclk21_i = '1') then
            tile0_tx_resetdone1_r  <= tile0_resetdone1_i   after DLY;
            tile0_tx_resetdone1_r2 <= tile0_tx_resetdone1_r   after DLY;
        end if;
    end process;

    



    ------------------------------ Frame Generators ---------------------------
    -- The example design uses Block RAM based frame generators to provide test
    -- data to the GTXs for transmission. By default the frame generators are 
    -- loaded with an incrementing data sequence that includes commas/alignment
    -- characters for alignment. If your protocol uses channel bonding, the 
    -- frame generator will also be preloaded with a channel bonding sequence.
    
    -- You can modify the data transmitted by changing the INIT values of the frame
    -- generator in this file. Pay careful attention to bit order and the spacing
    -- of your control and alignment characters.

    tile0_frame_gen1 : FRAME_GEN
    generic map
    (
        WORDS_IN_BRAM                   =>      EXAMPLE_WORDS_IN_BRAM,
        MEM_00                  =>  x"0000000600000005000000040000000300000002000000bc0000000100000000",
        MEM_01                  =>  x"0000000e0000000d0000000c0000000b0000000a000000090000000800000007",
        MEM_02                  =>  x"000000160000001500000014000000130000001200000011000000100000000f",
        MEM_03                  =>  x"0000001e0000001d0000001c0000001b0000001a000000190000001800000017",
        MEM_04                  =>  x"000000260000002500000024000000230000002200000021000000200000001f",
        MEM_05                  =>  x"0000002e0000002d0000002c0000002b0000002a000000290000002800000027",
        MEM_06                  =>  x"000000360000003500000034000000330000003200000031000000300000002f",
        MEM_07                  =>  x"0000003e0000003d0000003c0000003b0000003a000000390000003800000037",
        MEM_08                  =>  x"000000460000004500000044000000430000004200000041000000400000003f",
        MEM_09                  =>  x"0000004e0000004d0000004c0000004b0000004a000000490000004800000047",
        MEM_0A                  =>  x"000000560000005500000054000000530000005200000051000000500000004f",
        MEM_0B                  =>  x"0000005e0000005d0000005c0000005b0000005a000000590000005800000057",
        MEM_0C                  =>  x"000000660000006500000064000000630000006200000061000000600000005f",
        MEM_0D                  =>  x"0000006e0000006d0000006c0000006b0000006a000000690000006800000067",
        MEM_0E                  =>  x"000000760000007500000074000000730000007200000071000000700000006f",
        MEM_0F                  =>  x"0000007e0000007d0000007c0000007b0000007a000000790000007800000077",
        MEM_10                  =>  x"0000000600000005000000040000000300000002000000bc0000000100000000",
        MEM_11                  =>  x"0000000e0000000d0000000c0000000b0000000a000000090000000800000007",
        MEM_12                  =>  x"000000160000001500000014000000130000001200000011000000100000000f",
        MEM_13                  =>  x"0000001e0000001d0000001c0000001b0000001a000000190000001800000017",
        MEM_14                  =>  x"000000260000002500000024000000230000002200000021000000200000001f",
        MEM_15                  =>  x"0000002e0000002d0000002c0000002b0000002a000000290000002800000027",
        MEM_16                  =>  x"000000360000003500000034000000330000003200000031000000300000002f",
        MEM_17                  =>  x"0000003e0000003d0000003c0000003b0000003a000000390000003800000037",
        MEM_18                  =>  x"000000460000004500000044000000430000004200000041000000400000003f",
        MEM_19                  =>  x"0000004e0000004d0000004c0000004b0000004a000000490000004800000047",
        MEM_1A                  =>  x"000000560000005500000054000000530000005200000051000000500000004f",
        MEM_1B                  =>  x"0000005e0000005d0000005c0000005b0000005a000000590000005800000057",
        MEM_1C                  =>  x"000000660000006500000064000000630000006200000061000000600000005f",
        MEM_1D                  =>  x"0000006e0000006d0000006c0000006b0000006a000000690000006800000067",
        MEM_1E                  =>  x"000000760000007500000074000000730000007200000071000000700000006f",
        MEM_1F                  =>  x"0000007e0000007d0000007c0000007b0000007a000000790000007800000077",
        MEM_20                  =>  x"0000000600000005000000040000000300000002000000bc0000000100000000",
        MEM_21                  =>  x"0000000e0000000d0000000c0000000b0000000a000000090000000800000007",
        MEM_22                  =>  x"000000160000001500000014000000130000001200000011000000100000000f",
        MEM_23                  =>  x"0000001e0000001d0000001c0000001b0000001a000000190000001800000017",
        MEM_24                  =>  x"000000260000002500000024000000230000002200000021000000200000001f",
        MEM_25                  =>  x"0000002e0000002d0000002c0000002b0000002a000000290000002800000027",
        MEM_26                  =>  x"000000360000003500000034000000330000003200000031000000300000002f",
        MEM_27                  =>  x"0000003e0000003d0000003c0000003b0000003a000000390000003800000037",
        MEM_28                  =>  x"000000460000004500000044000000430000004200000041000000400000003f",
        MEM_29                  =>  x"0000004e0000004d0000004c0000004b0000004a000000490000004800000047",
        MEM_2A                  =>  x"000000560000005500000054000000530000005200000051000000500000004f",
        MEM_2B                  =>  x"0000005e0000005d0000005c0000005b0000005a000000590000005800000057",
        MEM_2C                  =>  x"000000660000006500000064000000630000006200000061000000600000005f",
        MEM_2D                  =>  x"0000006e0000006d0000006c0000006b0000006a000000690000006800000067",
        MEM_2E                  =>  x"000000760000007500000074000000730000007200000071000000700000006f",
        MEM_2F                  =>  x"0000007e0000007d0000007c0000007b0000007a000000790000007800000077",
        MEM_30                  =>  x"0000000600000005000000040000000300000002000000bc0000000100000000",
        MEM_31                  =>  x"0000000e0000000d0000000c0000000b0000000a000000090000000800000007",
        MEM_32                  =>  x"000000160000001500000014000000130000001200000011000000100000000f",
        MEM_33                  =>  x"0000001e0000001d0000001c0000001b0000001a000000190000001800000017",
        MEM_34                  =>  x"000000260000002500000024000000230000002200000021000000200000001f",
        MEM_35                  =>  x"0000002e0000002d0000002c0000002b0000002a000000290000002800000027",
        MEM_36                  =>  x"000000360000003500000034000000330000003200000031000000300000002f",
        MEM_37                  =>  x"0000003e0000003d0000003c0000003b0000003a000000390000003800000037",
        MEM_38                  =>  x"000000460000004500000044000000430000004200000041000000400000003f",
        MEM_39                  =>  x"0000004e0000004d0000004c0000004b0000004a000000490000004800000047",
        MEM_3A                  =>  x"000000560000005500000054000000530000005200000051000000500000004f",
        MEM_3B                  =>  x"0000005e0000005d0000005c0000005b0000005a000000590000005800000057",
        MEM_3C                  =>  x"000000660000006500000064000000630000006200000061000000600000005f",
        MEM_3D                  =>  x"0000006e0000006d0000006c0000006b0000006a000000690000006800000067",
        MEM_3E                  =>  x"000000760000007500000074000000730000007200000071000000700000006f",
        MEM_3F                  =>  x"0000007e0000007d0000007c0000007b0000007a000000790000007800000077",
        MEMP_00                  =>  x"0000000000000000000000000000000000000000000000000000000000000100",
        MEMP_01                  =>  x"0000000000000000000000000000000000000000000000000000000000000000",
        MEMP_02                  =>  x"0000000000000000000000000000000000000000000000000000000000000100",
        MEMP_03                  =>  x"0000000000000000000000000000000000000000000000000000000000000000",
        MEMP_04                  =>  x"0000000000000000000000000000000000000000000000000000000000000100",
        MEMP_05                  =>  x"0000000000000000000000000000000000000000000000000000000000000000",
        MEMP_06                  =>  x"0000000000000000000000000000000000000000000000000000000000000100",
        MEMP_07                  =>  x"0000000000000000000000000000000000000000000000000000000000000000"
    )
    port map
    (
        -- User Interface
        TX_DATA(39 downto 8)            =>      tile0_txdata1_float_i,
        TX_DATA(7 downto 0)             =>      tile0_txdata1_i,
 
        TX_CHARISK(3 downto 1)          =>      tile0_txcharisk1_float_i,
        TX_CHARISK(0)                   =>      tile0_txcharisk1_i,
        -- System Interface
        USER_CLK                        =>      tile0_txusrclk21_i,
        SYSTEM_RESET                    =>      tile0_tx_system_reset1_c
    );
    


    ---------------------------------- Frame Checkers -------------------------
    -- The example design uses Block RAM based frame checkers to verify incoming  
    -- data. By default the frame generators are loaded with a data sequence that 
    -- matches the outgoing sequence of the frame generators for the TX ports.
    
    -- You can modify the expected data sequence by changing the INIT values of the frame
    -- checkers in this file. Pay careful attention to bit order and the spacing
    -- of your control and alignment characters.
    
    -- When the frame checker receives data, it attempts to synchronise to the 
    -- incoming pattern by looking for the first sequence in the pattern. Once it 
    -- finds the first sequence, it increments through the sequence, and indicates an 
    -- error whenever the next value received does not match the expected value.

     -- This GTX is not active.The match port for pattern checker of this GTX is tied off
    tile0_matchn0_i                         <= '0';

    tile0_frame_check1_reset_i              <= reset_on_data_error_i when (EXAMPLE_CONFIG_INDEPENDENT_LANES=0) else tile0_matchn1_i;

    -- tile0_frame_check0 is always connected to the lane with the start of char
    -- and this lane starts off the data checking on all the other lanes. The INC_IN port is tied off
    tile0_inc_in1_i                         <= '0';

    tile0_frame_check1 : FRAME_CHECK
    generic map
    (
        RX_DATA_WIDTH                   =>      8,
        USE_COMMA                       =>      1,
        WORDS_IN_BRAM                   =>      EXAMPLE_WORDS_IN_BRAM,
        CONFIG_INDEPENDENT_LANES        =>      1,
        START_OF_PACKET_CHAR            =>      x"bc",
        MEM_00                  =>  x"0000000600000005000000040000000300000002000000bc0000000100000000",
        MEM_01                  =>  x"0000000e0000000d0000000c0000000b0000000a000000090000000800000007",
        MEM_02                  =>  x"000000160000001500000014000000130000001200000011000000100000000f",
        MEM_03                  =>  x"0000001e0000001d0000001c0000001b0000001a000000190000001800000017",
        MEM_04                  =>  x"000000260000002500000024000000230000002200000021000000200000001f",
        MEM_05                  =>  x"0000002e0000002d0000002c0000002b0000002a000000290000002800000027",
        MEM_06                  =>  x"000000360000003500000034000000330000003200000031000000300000002f",
        MEM_07                  =>  x"0000003e0000003d0000003c0000003b0000003a000000390000003800000037",
        MEM_08                  =>  x"000000460000004500000044000000430000004200000041000000400000003f",
        MEM_09                  =>  x"0000004e0000004d0000004c0000004b0000004a000000490000004800000047",
        MEM_0A                  =>  x"000000560000005500000054000000530000005200000051000000500000004f",
        MEM_0B                  =>  x"0000005e0000005d0000005c0000005b0000005a000000590000005800000057",
        MEM_0C                  =>  x"000000660000006500000064000000630000006200000061000000600000005f",
        MEM_0D                  =>  x"0000006e0000006d0000006c0000006b0000006a000000690000006800000067",
        MEM_0E                  =>  x"000000760000007500000074000000730000007200000071000000700000006f",
        MEM_0F                  =>  x"0000007e0000007d0000007c0000007b0000007a000000790000007800000077",
        MEM_10                  =>  x"0000000600000005000000040000000300000002000000bc0000000100000000",
        MEM_11                  =>  x"0000000e0000000d0000000c0000000b0000000a000000090000000800000007",
        MEM_12                  =>  x"000000160000001500000014000000130000001200000011000000100000000f",
        MEM_13                  =>  x"0000001e0000001d0000001c0000001b0000001a000000190000001800000017",
        MEM_14                  =>  x"000000260000002500000024000000230000002200000021000000200000001f",
        MEM_15                  =>  x"0000002e0000002d0000002c0000002b0000002a000000290000002800000027",
        MEM_16                  =>  x"000000360000003500000034000000330000003200000031000000300000002f",
        MEM_17                  =>  x"0000003e0000003d0000003c0000003b0000003a000000390000003800000037",
        MEM_18                  =>  x"000000460000004500000044000000430000004200000041000000400000003f",
        MEM_19                  =>  x"0000004e0000004d0000004c0000004b0000004a000000490000004800000047",
        MEM_1A                  =>  x"000000560000005500000054000000530000005200000051000000500000004f",
        MEM_1B                  =>  x"0000005e0000005d0000005c0000005b0000005a000000590000005800000057",
        MEM_1C                  =>  x"000000660000006500000064000000630000006200000061000000600000005f",
        MEM_1D                  =>  x"0000006e0000006d0000006c0000006b0000006a000000690000006800000067",
        MEM_1E                  =>  x"000000760000007500000074000000730000007200000071000000700000006f",
        MEM_1F                  =>  x"0000007e0000007d0000007c0000007b0000007a000000790000007800000077",
        MEM_20                  =>  x"0000000600000005000000040000000300000002000000bc0000000100000000",
        MEM_21                  =>  x"0000000e0000000d0000000c0000000b0000000a000000090000000800000007",
        MEM_22                  =>  x"000000160000001500000014000000130000001200000011000000100000000f",
        MEM_23                  =>  x"0000001e0000001d0000001c0000001b0000001a000000190000001800000017",
        MEM_24                  =>  x"000000260000002500000024000000230000002200000021000000200000001f",
        MEM_25                  =>  x"0000002e0000002d0000002c0000002b0000002a000000290000002800000027",
        MEM_26                  =>  x"000000360000003500000034000000330000003200000031000000300000002f",
        MEM_27                  =>  x"0000003e0000003d0000003c0000003b0000003a000000390000003800000037",
        MEM_28                  =>  x"000000460000004500000044000000430000004200000041000000400000003f",
        MEM_29                  =>  x"0000004e0000004d0000004c0000004b0000004a000000490000004800000047",
        MEM_2A                  =>  x"000000560000005500000054000000530000005200000051000000500000004f",
        MEM_2B                  =>  x"0000005e0000005d0000005c0000005b0000005a000000590000005800000057",
        MEM_2C                  =>  x"000000660000006500000064000000630000006200000061000000600000005f",
        MEM_2D                  =>  x"0000006e0000006d0000006c0000006b0000006a000000690000006800000067",
        MEM_2E                  =>  x"000000760000007500000074000000730000007200000071000000700000006f",
        MEM_2F                  =>  x"0000007e0000007d0000007c0000007b0000007a000000790000007800000077",
        MEM_30                  =>  x"0000000600000005000000040000000300000002000000bc0000000100000000",
        MEM_31                  =>  x"0000000e0000000d0000000c0000000b0000000a000000090000000800000007",
        MEM_32                  =>  x"000000160000001500000014000000130000001200000011000000100000000f",
        MEM_33                  =>  x"0000001e0000001d0000001c0000001b0000001a000000190000001800000017",
        MEM_34                  =>  x"000000260000002500000024000000230000002200000021000000200000001f",
        MEM_35                  =>  x"0000002e0000002d0000002c0000002b0000002a000000290000002800000027",
        MEM_36                  =>  x"000000360000003500000034000000330000003200000031000000300000002f",
        MEM_37                  =>  x"0000003e0000003d0000003c0000003b0000003a000000390000003800000037",
        MEM_38                  =>  x"000000460000004500000044000000430000004200000041000000400000003f",
        MEM_39                  =>  x"0000004e0000004d0000004c0000004b0000004a000000490000004800000047",
        MEM_3A                  =>  x"000000560000005500000054000000530000005200000051000000500000004f",
        MEM_3B                  =>  x"0000005e0000005d0000005c0000005b0000005a000000590000005800000057",
        MEM_3C                  =>  x"000000660000006500000064000000630000006200000061000000600000005f",
        MEM_3D                  =>  x"0000006e0000006d0000006c0000006b0000006a000000690000006800000067",
        MEM_3E                  =>  x"000000760000007500000074000000730000007200000071000000700000006f",
        MEM_3F                  =>  x"0000007e0000007d0000007c0000007b0000007a000000790000007800000077",
        MEMP_00                  =>  x"0000000000000000000000000000000000000000000000000000000000000100",
        MEMP_01                  =>  x"0000000000000000000000000000000000000000000000000000000000000000",
        MEMP_02                  =>  x"0000000000000000000000000000000000000000000000000000000000000100",
        MEMP_03                  =>  x"0000000000000000000000000000000000000000000000000000000000000000",
        MEMP_04                  =>  x"0000000000000000000000000000000000000000000000000000000000000100",
        MEMP_05                  =>  x"0000000000000000000000000000000000000000000000000000000000000000",
        MEMP_06                  =>  x"0000000000000000000000000000000000000000000000000000000000000100",
        MEMP_07                  =>  x"0000000000000000000000000000000000000000000000000000000000000000"
    )
    port map
    (
        -- MGT Interface
        RX_DATA                         =>      tile0_rxdata1_i,
        RX_ENMCOMMA_ALIGN               =>      tile0_rxenmcommaalign1_i,
        RX_ENPCOMMA_ALIGN               =>      tile0_rxenpcommaalign1_i,
        RX_ENCHAN_SYNC                  =>      open,
        RX_CHANBOND_SEQ                 =>      tied_to_ground_i,
        -- Control Interface
        INC_IN                          =>      tile0_inc_in1_i,
        INC_OUT                         =>      tile0_inc_out1_i,
        PATTERN_MATCH_N                 =>      tile0_matchn1_i,
        RESET_ON_ERROR                  =>      tile0_frame_check1_reset_i,
        -- System Interface
        USER_CLK                        =>      tile0_txusrclk21_i,
        SYSTEM_RESET                    =>      tile0_rx_system_reset1_c,
        ERROR_COUNT                     =>      tile0_error_count1_i
    );
        





    ----------------------------- Chipscope Connections -----------------------
    -- When the example design is run in hardware, it uses chipscope to allow the
    -- example design and GTX wrapper to be controlled and monitored. The 
    -- EXAMPLE_USE_CHIPSCOPE parameter allows chipscope to be removed for simulation.
    
chipscope : if EXAMPLE_USE_CHIPSCOPE = 1 generate


    -- Shared VIO for all tiles
    shared_vio_i : shared_vio
    port map
    (
        control                         =>      shared_vio_control_i,
        async_in                        =>      shared_vio_in_i,
        async_out                       =>      shared_vio_out_i
    );

    -- ICON for all VIOs 
    i_icon : icon
    port map
    (
        control0                        =>      shared_vio_control_i,
        control1                        =>      tx_data_vio_control0_i,
        control2                        =>      rx_data_vio_control0_i,
        control3                        =>      ila_control0_i,
        control4                        =>      tx_data_vio_control1_i,
        control5                        =>      rx_data_vio_control1_i,
        control6                        =>      ila_control1_i
    );

    -- TX VIO 
    tx_data_vio0_i : shared_vio
    port map
    (
        control                         =>      tx_data_vio_control0_i,
        async_in                        =>      tx_data_vio_in0_i,
        async_out                       =>      tx_data_vio_out0_i
    );
    
    -- RX VIO 
    rx_data_vio0_i : shared_vio
    port map
    (
        control                         =>      rx_data_vio_control0_i,
        async_in                        =>      rx_data_vio_in0_i,
        async_out                       =>      rx_data_vio_out0_i
    );
    
    -- RX ILA
    ila0_i : ila
    port map
    (
        control                         =>      ila_control0_i,
        clk                             =>      ila_clk0_i,
        trig0                           =>      ila_in0_i
    );

    
    -- The RX ILA must use the same clock as the selected transceiver
    ila_clk0_bufg_i : BUFG
    port map
    (
        I => ila_clk_mux_out0_i,
        O => ila_clk0_i
    );

     ila_clk_mux_out0_i <= '0';


    -- TX VIO 
    tx_data_vio1_i : shared_vio
    port map
    (
        control                         =>      tx_data_vio_control1_i,
        async_in                        =>      tx_data_vio_in1_i,
        async_out                       =>      tx_data_vio_out1_i
    );
    
    -- RX VIO 
    rx_data_vio1_i : shared_vio
    port map
    (
        control                         =>      rx_data_vio_control1_i,
        async_in                        =>      rx_data_vio_in1_i,
        async_out                       =>      rx_data_vio_out1_i
    );
    
    -- RX ILA
    ila1_i : ila
    port map
    (
        control                         =>      ila_control1_i,
        clk                             =>      ila_clk1_i,
        trig0                           =>      ila_in1_i
    );

    
    -- The RX ILA must use the same clock as the selected transceiver
    ila_clk1_bufg_i : BUFG
    port map
    (
        I => ila_clk_mux_out1_i,
        O => ila_clk1_i
    );

     ila_clk_mux_out1_i <= tile0_txusrclk21_i;



    -- assign resets for frame_gen modules
    tile0_tx_system_reset1_c                <= not tile0_tx_resetdone1_r2 or user_tx_reset_i;
    -- assign resets for frame_check modules
    tile0_rx_system_reset1_c                <= not tile0_rx_resetdone1_r2 or user_rx_reset_i;


    tile0_gtxreset_i                        <= gtxreset_i;

    -- Shared VIO Outputs
    gtxreset_i                              <= shared_vio_out_i(31);
    user_tx_reset_i                         <= shared_vio_out_i(30);
    user_rx_reset_i                         <= shared_vio_out_i(29);

    -- Shared VIO Inputs
    shared_vio_in_i(31)                     <= tile0_plllkdet_i;
    shared_vio_in_i(30 downto 0)            <= "0000000000000000000000000000000";

    -- Chipscope connections for GTP0 on Tile 0
    tile0_tx_data_vio_in0_i(31 downto 0)    <= "00000000000000000000000000000000";
    tile0_loopback0_i                       <= tx_data_vio_out0_i(31 downto 29);
    tile0_rx_data_vio_in0_i(31)             <= tile0_resetdone0_i;
    tile0_rx_data_vio_in0_i(30 downto 0)    <= "0000000000000000000000000000000";
    tile0_ila_in0_i(84 downto 77)           <= tile0_error_count0_i;
    tile0_ila_in0_i(76 downto 0)            <= "00000000000000000000000000000000000000000000000000000000000000000000000000000";

    -- Chipscope connections for GTP1 on Tile 0
    tile0_tx_data_vio_in1_i(31 downto 0)    <= "00000000000000000000000000000000";
    tile0_loopback1_i                       <= tx_data_vio_out1_i(31 downto 29);
    tile0_rx_data_vio_in1_i(31)             <= tile0_resetdone1_i;
    tile0_rx_data_vio_in1_i(30 downto 0)    <= "0000000000000000000000000000000";
    tile0_ila_in1_i(84)                     <= tile0_rxcharisk1_i;
    tile0_ila_in1_i(83)                     <= tile0_rxdisperr1_i;
    tile0_ila_in1_i(82)                     <= tile0_rxnotintable1_i;
    tile0_ila_in1_i(81 downto 79)           <= tile0_rxclkcorcnt1_i;
    tile0_ila_in1_i(78 downto 71)           <= tile0_rxdata1_i;
    tile0_ila_in1_i(70 downto 69)           <= tile0_rxlossofsync1_i;
    tile0_ila_in1_i(68 downto 61)           <= tile0_error_count1_i;
    tile0_ila_in1_i(60 downto 0)            <= "0000000000000000000000000000000000000000000000000000000000000";


    tx_data_vio_in0_i                   <=      tile0_tx_data_vio_in0_i;


    rx_data_vio_in0_i                   <=      tile0_rx_data_vio_in0_i;


    ila_in0_i                           <=      tile0_ila_in0_i;



    tx_data_vio_in1_i                   <=      tile0_tx_data_vio_in1_i;


    rx_data_vio_in1_i                   <=      tile0_rx_data_vio_in1_i;


    ila_in1_i                           <=      tile0_ila_in1_i;





   
end generate chipscope;


no_chipscope : if EXAMPLE_USE_CHIPSCOPE = 0 generate

    -- If Chipscope is not being used, drive GTX reset signal
    -- from the top level ports
    tile0_gtxreset_i                        <= GTXRESET_IN;

    -- assign resets for frame_gen modules
    tile0_tx_system_reset1_c                <= not tile0_tx_resetdone1_r2;
    -- assign resets for frame_check modules
    tile0_rx_system_reset1_c                <= not tile0_rx_resetdone1_r2;

    gtxreset_i                              <= tied_to_ground_i;
    user_tx_reset_i                         <= tied_to_ground_i;
    user_rx_reset_i                         <= tied_to_ground_i;
    tile0_loopback0_i                       <= tied_to_ground_vec_i(2 downto 0);
    tile0_loopback1_i                       <= tied_to_ground_vec_i(2 downto 0);



end generate no_chipscope;


end RTL;


