------------------------------------------------------------------------------_
--$Date: 2008/05/30 00:57:53 $
--$RCSfile: mgt_usrclk_source_dcm_vhd.ejava,v $
--$Revision: 1.1.2.1 $
-------------------------------------------------------------------------------
--   __  __ 
--  /   /\/   / 
-- /__/  \   /    Vendor: Xilinx 
-- \   \   \/     Version : 1.5
--  \   \         Application : RocketIO GTX Wizard 
--  /   /         Filename : mgt_usrclk_source.vhd
-- /__/   /\      Timestamp : 02/08/2005 09:12:43
-- \   \  /  \ 
--  \__\/\__\ 
--
--
-- Module MGT_USRCLK_SOURCE (for use with GTX Transceivers)
-- Generated by Xilinx RocketIO GTX Wizard

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;


--***********************************Entity Declaration************************
entity MGT_USRCLK_SOURCE is
generic
(
    FREQUENCY_MODE     : string   := "LOW";    
    PERFORMANCE_MODE   : string   := "MAX_SPEED"    
);
port
(
    DIV1_OUT                : out std_logic;
    DIV2_OUT                : out std_logic;
    DCM_LOCKED_OUT          : out std_logic;
    CLK_IN                  : in  std_logic;
    DCM_RESET_IN            : in  std_logic

);

    attribute X_CORE_INFO : string;
    attribute X_CORE_INFO of MGT_USRCLK_SOURCE : entity is "gtxwizard_v1_5, Coregen v10.1_ip3";

end MGT_USRCLK_SOURCE;

architecture RTL of MGT_USRCLK_SOURCE is
--*********************************Wire Declarations***************************

    signal not_connected_i          : std_logic_vector(15 downto 0);
    signal clkfb_i                  : std_logic;
    signal clkdv_i                  : std_logic;
    signal clk0_i                   : std_logic;
    signal tied_to_ground_i         : std_logic;
    signal tied_to_ground_vec_i     : std_logic_vector(63 downto 0);

begin

--*********************************** Main Body of Code ***********************


    --  Static signal Assigments    
    tied_to_ground_i                  <= '0';        
    tied_to_ground_vec_i(63 downto 0) <= (others => '0');

    -- Instantiate a DCM module to divide the reference clock.
    clock_divider_i : DCM_BASE
    generic map
    (
        CLKDV_DIVIDE          =>          2.0,
        DFS_FREQUENCY_MODE    =>          "LOW", 
        DLL_FREQUENCY_MODE    =>          FREQUENCY_MODE,
        DCM_PERFORMANCE_MODE  =>          PERFORMANCE_MODE
    )    
    port map
    (
        CLK0                =>          clk0_i,
        CLK180              =>          open,
        CLK270              =>          open,
        CLK2X               =>          open,
        CLK2X180            =>          open,
        CLK90               =>          open,
        CLKDV               =>          clkdv_i,
        CLKFX               =>          open,
        CLKFX180            =>          open,
        LOCKED              =>          DCM_LOCKED_OUT,
        CLKFB               =>          clkfb_i,
        CLKIN               =>          CLK_IN,
        RST                 =>          DCM_RESET_IN
    );


    dcm_1x_bufg_i : BUFG
    port map
    (
        I                   =>          clk0_i,
        O                   =>          clkfb_i
    );
    
    
    DIV1_OUT  <=  clkfb_i;


    dcm_div2_bufg_i : BUFG 
    port map
    (
        I                   =>          clkdv_i,
        O                   =>          DIV2_OUT
    );



end RTL;

